module GenTanh(
	input [15:0] x,
	output reg [15:0] y
);

	always @(*) begin
		case(x)
			16'h8000: y = 16'hfe00;
			16'h8001: y = 16'hfe00;
			16'h8002: y = 16'hfe00;
			16'h8003: y = 16'hfe00;
			16'h8004: y = 16'hfe00;
			16'h8005: y = 16'hfe00;
			16'h8006: y = 16'hfe00;
			16'h8007: y = 16'hfe00;
			16'h8008: y = 16'hfe00;
			16'h8009: y = 16'hfe00;
			16'h800a: y = 16'hfe00;
			16'h800b: y = 16'hfe00;
			16'h800c: y = 16'hfe00;
			16'h800d: y = 16'hfe00;
			16'h800e: y = 16'hfe00;
			16'h800f: y = 16'hfe00;
			16'h8010: y = 16'hfe00;
			16'h8011: y = 16'hfe00;
			16'h8012: y = 16'hfe00;
			16'h8013: y = 16'hfe00;
			16'h8014: y = 16'hfe00;
			16'h8015: y = 16'hfe00;
			16'h8016: y = 16'hfe00;
			16'h8017: y = 16'hfe00;
			16'h8018: y = 16'hfe00;
			16'h8019: y = 16'hfe00;
			16'h801a: y = 16'hfe00;
			16'h801b: y = 16'hfe00;
			16'h801c: y = 16'hfe00;
			16'h801d: y = 16'hfe00;
			16'h801e: y = 16'hfe00;
			16'h801f: y = 16'hfe00;
			16'h8020: y = 16'hfe00;
			16'h8021: y = 16'hfe00;
			16'h8022: y = 16'hfe00;
			16'h8023: y = 16'hfe00;
			16'h8024: y = 16'hfe00;
			16'h8025: y = 16'hfe00;
			16'h8026: y = 16'hfe00;
			16'h8027: y = 16'hfe00;
			16'h8028: y = 16'hfe00;
			16'h8029: y = 16'hfe00;
			16'h802a: y = 16'hfe00;
			16'h802b: y = 16'hfe00;
			16'h802c: y = 16'hfe00;
			16'h802d: y = 16'hfe00;
			16'h802e: y = 16'hfe00;
			16'h802f: y = 16'hfe00;
			16'h8030: y = 16'hfe00;
			16'h8031: y = 16'hfe00;
			16'h8032: y = 16'hfe00;
			16'h8033: y = 16'hfe00;
			16'h8034: y = 16'hfe00;
			16'h8035: y = 16'hfe00;
			16'h8036: y = 16'hfe00;
			16'h8037: y = 16'hfe00;
			16'h8038: y = 16'hfe00;
			16'h8039: y = 16'hfe00;
			16'h803a: y = 16'hfe00;
			16'h803b: y = 16'hfe00;
			16'h803c: y = 16'hfe00;
			16'h803d: y = 16'hfe00;
			16'h803e: y = 16'hfe00;
			16'h803f: y = 16'hfe00;
			16'h8040: y = 16'hfe00;
			16'h8041: y = 16'hfe00;
			16'h8042: y = 16'hfe00;
			16'h8043: y = 16'hfe00;
			16'h8044: y = 16'hfe00;
			16'h8045: y = 16'hfe00;
			16'h8046: y = 16'hfe00;
			16'h8047: y = 16'hfe00;
			16'h8048: y = 16'hfe00;
			16'h8049: y = 16'hfe00;
			16'h804a: y = 16'hfe00;
			16'h804b: y = 16'hfe00;
			16'h804c: y = 16'hfe00;
			16'h804d: y = 16'hfe00;
			16'h804e: y = 16'hfe00;
			16'h804f: y = 16'hfe00;
			16'h8050: y = 16'hfe00;
			16'h8051: y = 16'hfe00;
			16'h8052: y = 16'hfe00;
			16'h8053: y = 16'hfe00;
			16'h8054: y = 16'hfe00;
			16'h8055: y = 16'hfe00;
			16'h8056: y = 16'hfe00;
			16'h8057: y = 16'hfe00;
			16'h8058: y = 16'hfe00;
			16'h8059: y = 16'hfe00;
			16'h805a: y = 16'hfe00;
			16'h805b: y = 16'hfe00;
			16'h805c: y = 16'hfe00;
			16'h805d: y = 16'hfe00;
			16'h805e: y = 16'hfe00;
			16'h805f: y = 16'hfe00;
			16'h8060: y = 16'hfe00;
			16'h8061: y = 16'hfe00;
			16'h8062: y = 16'hfe00;
			16'h8063: y = 16'hfe00;
			16'h8064: y = 16'hfe00;
			16'h8065: y = 16'hfe00;
			16'h8066: y = 16'hfe00;
			16'h8067: y = 16'hfe00;
			16'h8068: y = 16'hfe00;
			16'h8069: y = 16'hfe00;
			16'h806a: y = 16'hfe00;
			16'h806b: y = 16'hfe00;
			16'h806c: y = 16'hfe00;
			16'h806d: y = 16'hfe00;
			16'h806e: y = 16'hfe00;
			16'h806f: y = 16'hfe00;
			16'h8070: y = 16'hfe00;
			16'h8071: y = 16'hfe00;
			16'h8072: y = 16'hfe00;
			16'h8073: y = 16'hfe00;
			16'h8074: y = 16'hfe00;
			16'h8075: y = 16'hfe00;
			16'h8076: y = 16'hfe00;
			16'h8077: y = 16'hfe00;
			16'h8078: y = 16'hfe00;
			16'h8079: y = 16'hfe00;
			16'h807a: y = 16'hfe00;
			16'h807b: y = 16'hfe00;
			16'h807c: y = 16'hfe00;
			16'h807d: y = 16'hfe00;
			16'h807e: y = 16'hfe00;
			16'h807f: y = 16'hfe00;
			16'h8080: y = 16'hfe00;
			16'h8081: y = 16'hfe00;
			16'h8082: y = 16'hfe00;
			16'h8083: y = 16'hfe00;
			16'h8084: y = 16'hfe00;
			16'h8085: y = 16'hfe00;
			16'h8086: y = 16'hfe00;
			16'h8087: y = 16'hfe00;
			16'h8088: y = 16'hfe00;
			16'h8089: y = 16'hfe00;
			16'h808a: y = 16'hfe00;
			16'h808b: y = 16'hfe00;
			16'h808c: y = 16'hfe00;
			16'h808d: y = 16'hfe00;
			16'h808e: y = 16'hfe00;
			16'h808f: y = 16'hfe00;
			16'h8090: y = 16'hfe00;
			16'h8091: y = 16'hfe00;
			16'h8092: y = 16'hfe00;
			16'h8093: y = 16'hfe00;
			16'h8094: y = 16'hfe00;
			16'h8095: y = 16'hfe00;
			16'h8096: y = 16'hfe00;
			16'h8097: y = 16'hfe00;
			16'h8098: y = 16'hfe00;
			16'h8099: y = 16'hfe00;
			16'h809a: y = 16'hfe00;
			16'h809b: y = 16'hfe00;
			16'h809c: y = 16'hfe00;
			16'h809d: y = 16'hfe00;
			16'h809e: y = 16'hfe00;
			16'h809f: y = 16'hfe00;
			16'h80a0: y = 16'hfe00;
			16'h80a1: y = 16'hfe00;
			16'h80a2: y = 16'hfe00;
			16'h80a3: y = 16'hfe00;
			16'h80a4: y = 16'hfe00;
			16'h80a5: y = 16'hfe00;
			16'h80a6: y = 16'hfe00;
			16'h80a7: y = 16'hfe00;
			16'h80a8: y = 16'hfe00;
			16'h80a9: y = 16'hfe00;
			16'h80aa: y = 16'hfe00;
			16'h80ab: y = 16'hfe00;
			16'h80ac: y = 16'hfe00;
			16'h80ad: y = 16'hfe00;
			16'h80ae: y = 16'hfe00;
			16'h80af: y = 16'hfe00;
			16'h80b0: y = 16'hfe00;
			16'h80b1: y = 16'hfe00;
			16'h80b2: y = 16'hfe00;
			16'h80b3: y = 16'hfe00;
			16'h80b4: y = 16'hfe00;
			16'h80b5: y = 16'hfe00;
			16'h80b6: y = 16'hfe00;
			16'h80b7: y = 16'hfe00;
			16'h80b8: y = 16'hfe00;
			16'h80b9: y = 16'hfe00;
			16'h80ba: y = 16'hfe00;
			16'h80bb: y = 16'hfe00;
			16'h80bc: y = 16'hfe00;
			16'h80bd: y = 16'hfe00;
			16'h80be: y = 16'hfe00;
			16'h80bf: y = 16'hfe00;
			16'h80c0: y = 16'hfe00;
			16'h80c1: y = 16'hfe00;
			16'h80c2: y = 16'hfe00;
			16'h80c3: y = 16'hfe00;
			16'h80c4: y = 16'hfe00;
			16'h80c5: y = 16'hfe00;
			16'h80c6: y = 16'hfe00;
			16'h80c7: y = 16'hfe00;
			16'h80c8: y = 16'hfe00;
			16'h80c9: y = 16'hfe00;
			16'h80ca: y = 16'hfe00;
			16'h80cb: y = 16'hfe00;
			16'h80cc: y = 16'hfe00;
			16'h80cd: y = 16'hfe00;
			16'h80ce: y = 16'hfe00;
			16'h80cf: y = 16'hfe00;
			16'h80d0: y = 16'hfe00;
			16'h80d1: y = 16'hfe00;
			16'h80d2: y = 16'hfe00;
			16'h80d3: y = 16'hfe00;
			16'h80d4: y = 16'hfe00;
			16'h80d5: y = 16'hfe00;
			16'h80d6: y = 16'hfe00;
			16'h80d7: y = 16'hfe00;
			16'h80d8: y = 16'hfe00;
			16'h80d9: y = 16'hfe00;
			16'h80da: y = 16'hfe00;
			16'h80db: y = 16'hfe00;
			16'h80dc: y = 16'hfe00;
			16'h80dd: y = 16'hfe00;
			16'h80de: y = 16'hfe00;
			16'h80df: y = 16'hfe00;
			16'h80e0: y = 16'hfe00;
			16'h80e1: y = 16'hfe00;
			16'h80e2: y = 16'hfe00;
			16'h80e3: y = 16'hfe00;
			16'h80e4: y = 16'hfe00;
			16'h80e5: y = 16'hfe00;
			16'h80e6: y = 16'hfe00;
			16'h80e7: y = 16'hfe00;
			16'h80e8: y = 16'hfe00;
			16'h80e9: y = 16'hfe00;
			16'h80ea: y = 16'hfe00;
			16'h80eb: y = 16'hfe00;
			16'h80ec: y = 16'hfe00;
			16'h80ed: y = 16'hfe00;
			16'h80ee: y = 16'hfe00;
			16'h80ef: y = 16'hfe00;
			16'h80f0: y = 16'hfe00;
			16'h80f1: y = 16'hfe00;
			16'h80f2: y = 16'hfe00;
			16'h80f3: y = 16'hfe00;
			16'h80f4: y = 16'hfe00;
			16'h80f5: y = 16'hfe00;
			16'h80f6: y = 16'hfe00;
			16'h80f7: y = 16'hfe00;
			16'h80f8: y = 16'hfe00;
			16'h80f9: y = 16'hfe00;
			16'h80fa: y = 16'hfe00;
			16'h80fb: y = 16'hfe00;
			16'h80fc: y = 16'hfe00;
			16'h80fd: y = 16'hfe00;
			16'h80fe: y = 16'hfe00;
			16'h80ff: y = 16'hfe00;
			16'h8100: y = 16'hfe00;
			16'h8101: y = 16'hfe00;
			16'h8102: y = 16'hfe00;
			16'h8103: y = 16'hfe00;
			16'h8104: y = 16'hfe00;
			16'h8105: y = 16'hfe00;
			16'h8106: y = 16'hfe00;
			16'h8107: y = 16'hfe00;
			16'h8108: y = 16'hfe00;
			16'h8109: y = 16'hfe00;
			16'h810a: y = 16'hfe00;
			16'h810b: y = 16'hfe00;
			16'h810c: y = 16'hfe00;
			16'h810d: y = 16'hfe00;
			16'h810e: y = 16'hfe00;
			16'h810f: y = 16'hfe00;
			16'h8110: y = 16'hfe00;
			16'h8111: y = 16'hfe00;
			16'h8112: y = 16'hfe00;
			16'h8113: y = 16'hfe00;
			16'h8114: y = 16'hfe00;
			16'h8115: y = 16'hfe00;
			16'h8116: y = 16'hfe00;
			16'h8117: y = 16'hfe00;
			16'h8118: y = 16'hfe00;
			16'h8119: y = 16'hfe00;
			16'h811a: y = 16'hfe00;
			16'h811b: y = 16'hfe00;
			16'h811c: y = 16'hfe00;
			16'h811d: y = 16'hfe00;
			16'h811e: y = 16'hfe00;
			16'h811f: y = 16'hfe00;
			16'h8120: y = 16'hfe00;
			16'h8121: y = 16'hfe00;
			16'h8122: y = 16'hfe00;
			16'h8123: y = 16'hfe00;
			16'h8124: y = 16'hfe00;
			16'h8125: y = 16'hfe00;
			16'h8126: y = 16'hfe00;
			16'h8127: y = 16'hfe00;
			16'h8128: y = 16'hfe00;
			16'h8129: y = 16'hfe00;
			16'h812a: y = 16'hfe00;
			16'h812b: y = 16'hfe00;
			16'h812c: y = 16'hfe00;
			16'h812d: y = 16'hfe00;
			16'h812e: y = 16'hfe00;
			16'h812f: y = 16'hfe00;
			16'h8130: y = 16'hfe00;
			16'h8131: y = 16'hfe00;
			16'h8132: y = 16'hfe00;
			16'h8133: y = 16'hfe00;
			16'h8134: y = 16'hfe00;
			16'h8135: y = 16'hfe00;
			16'h8136: y = 16'hfe00;
			16'h8137: y = 16'hfe00;
			16'h8138: y = 16'hfe00;
			16'h8139: y = 16'hfe00;
			16'h813a: y = 16'hfe00;
			16'h813b: y = 16'hfe00;
			16'h813c: y = 16'hfe00;
			16'h813d: y = 16'hfe00;
			16'h813e: y = 16'hfe00;
			16'h813f: y = 16'hfe00;
			16'h8140: y = 16'hfe00;
			16'h8141: y = 16'hfe00;
			16'h8142: y = 16'hfe00;
			16'h8143: y = 16'hfe00;
			16'h8144: y = 16'hfe00;
			16'h8145: y = 16'hfe00;
			16'h8146: y = 16'hfe00;
			16'h8147: y = 16'hfe00;
			16'h8148: y = 16'hfe00;
			16'h8149: y = 16'hfe00;
			16'h814a: y = 16'hfe00;
			16'h814b: y = 16'hfe00;
			16'h814c: y = 16'hfe00;
			16'h814d: y = 16'hfe00;
			16'h814e: y = 16'hfe00;
			16'h814f: y = 16'hfe00;
			16'h8150: y = 16'hfe00;
			16'h8151: y = 16'hfe00;
			16'h8152: y = 16'hfe00;
			16'h8153: y = 16'hfe00;
			16'h8154: y = 16'hfe00;
			16'h8155: y = 16'hfe00;
			16'h8156: y = 16'hfe00;
			16'h8157: y = 16'hfe00;
			16'h8158: y = 16'hfe00;
			16'h8159: y = 16'hfe00;
			16'h815a: y = 16'hfe00;
			16'h815b: y = 16'hfe00;
			16'h815c: y = 16'hfe00;
			16'h815d: y = 16'hfe00;
			16'h815e: y = 16'hfe00;
			16'h815f: y = 16'hfe00;
			16'h8160: y = 16'hfe00;
			16'h8161: y = 16'hfe00;
			16'h8162: y = 16'hfe00;
			16'h8163: y = 16'hfe00;
			16'h8164: y = 16'hfe00;
			16'h8165: y = 16'hfe00;
			16'h8166: y = 16'hfe00;
			16'h8167: y = 16'hfe00;
			16'h8168: y = 16'hfe00;
			16'h8169: y = 16'hfe00;
			16'h816a: y = 16'hfe00;
			16'h816b: y = 16'hfe00;
			16'h816c: y = 16'hfe00;
			16'h816d: y = 16'hfe00;
			16'h816e: y = 16'hfe00;
			16'h816f: y = 16'hfe00;
			16'h8170: y = 16'hfe00;
			16'h8171: y = 16'hfe00;
			16'h8172: y = 16'hfe00;
			16'h8173: y = 16'hfe00;
			16'h8174: y = 16'hfe00;
			16'h8175: y = 16'hfe00;
			16'h8176: y = 16'hfe00;
			16'h8177: y = 16'hfe00;
			16'h8178: y = 16'hfe00;
			16'h8179: y = 16'hfe00;
			16'h817a: y = 16'hfe00;
			16'h817b: y = 16'hfe00;
			16'h817c: y = 16'hfe00;
			16'h817d: y = 16'hfe00;
			16'h817e: y = 16'hfe00;
			16'h817f: y = 16'hfe00;
			16'h8180: y = 16'hfe00;
			16'h8181: y = 16'hfe00;
			16'h8182: y = 16'hfe00;
			16'h8183: y = 16'hfe00;
			16'h8184: y = 16'hfe00;
			16'h8185: y = 16'hfe00;
			16'h8186: y = 16'hfe00;
			16'h8187: y = 16'hfe00;
			16'h8188: y = 16'hfe00;
			16'h8189: y = 16'hfe00;
			16'h818a: y = 16'hfe00;
			16'h818b: y = 16'hfe00;
			16'h818c: y = 16'hfe00;
			16'h818d: y = 16'hfe00;
			16'h818e: y = 16'hfe00;
			16'h818f: y = 16'hfe00;
			16'h8190: y = 16'hfe00;
			16'h8191: y = 16'hfe00;
			16'h8192: y = 16'hfe00;
			16'h8193: y = 16'hfe00;
			16'h8194: y = 16'hfe00;
			16'h8195: y = 16'hfe00;
			16'h8196: y = 16'hfe00;
			16'h8197: y = 16'hfe00;
			16'h8198: y = 16'hfe00;
			16'h8199: y = 16'hfe00;
			16'h819a: y = 16'hfe00;
			16'h819b: y = 16'hfe00;
			16'h819c: y = 16'hfe00;
			16'h819d: y = 16'hfe00;
			16'h819e: y = 16'hfe00;
			16'h819f: y = 16'hfe00;
			16'h81a0: y = 16'hfe00;
			16'h81a1: y = 16'hfe00;
			16'h81a2: y = 16'hfe00;
			16'h81a3: y = 16'hfe00;
			16'h81a4: y = 16'hfe00;
			16'h81a5: y = 16'hfe00;
			16'h81a6: y = 16'hfe00;
			16'h81a7: y = 16'hfe00;
			16'h81a8: y = 16'hfe00;
			16'h81a9: y = 16'hfe00;
			16'h81aa: y = 16'hfe00;
			16'h81ab: y = 16'hfe00;
			16'h81ac: y = 16'hfe00;
			16'h81ad: y = 16'hfe00;
			16'h81ae: y = 16'hfe00;
			16'h81af: y = 16'hfe00;
			16'h81b0: y = 16'hfe00;
			16'h81b1: y = 16'hfe00;
			16'h81b2: y = 16'hfe00;
			16'h81b3: y = 16'hfe00;
			16'h81b4: y = 16'hfe00;
			16'h81b5: y = 16'hfe00;
			16'h81b6: y = 16'hfe00;
			16'h81b7: y = 16'hfe00;
			16'h81b8: y = 16'hfe00;
			16'h81b9: y = 16'hfe00;
			16'h81ba: y = 16'hfe00;
			16'h81bb: y = 16'hfe00;
			16'h81bc: y = 16'hfe00;
			16'h81bd: y = 16'hfe00;
			16'h81be: y = 16'hfe00;
			16'h81bf: y = 16'hfe00;
			16'h81c0: y = 16'hfe00;
			16'h81c1: y = 16'hfe00;
			16'h81c2: y = 16'hfe00;
			16'h81c3: y = 16'hfe00;
			16'h81c4: y = 16'hfe00;
			16'h81c5: y = 16'hfe00;
			16'h81c6: y = 16'hfe00;
			16'h81c7: y = 16'hfe00;
			16'h81c8: y = 16'hfe00;
			16'h81c9: y = 16'hfe00;
			16'h81ca: y = 16'hfe00;
			16'h81cb: y = 16'hfe00;
			16'h81cc: y = 16'hfe00;
			16'h81cd: y = 16'hfe00;
			16'h81ce: y = 16'hfe00;
			16'h81cf: y = 16'hfe00;
			16'h81d0: y = 16'hfe00;
			16'h81d1: y = 16'hfe00;
			16'h81d2: y = 16'hfe00;
			16'h81d3: y = 16'hfe00;
			16'h81d4: y = 16'hfe00;
			16'h81d5: y = 16'hfe00;
			16'h81d6: y = 16'hfe00;
			16'h81d7: y = 16'hfe00;
			16'h81d8: y = 16'hfe00;
			16'h81d9: y = 16'hfe00;
			16'h81da: y = 16'hfe00;
			16'h81db: y = 16'hfe00;
			16'h81dc: y = 16'hfe00;
			16'h81dd: y = 16'hfe00;
			16'h81de: y = 16'hfe00;
			16'h81df: y = 16'hfe00;
			16'h81e0: y = 16'hfe00;
			16'h81e1: y = 16'hfe00;
			16'h81e2: y = 16'hfe00;
			16'h81e3: y = 16'hfe00;
			16'h81e4: y = 16'hfe00;
			16'h81e5: y = 16'hfe00;
			16'h81e6: y = 16'hfe00;
			16'h81e7: y = 16'hfe00;
			16'h81e8: y = 16'hfe00;
			16'h81e9: y = 16'hfe00;
			16'h81ea: y = 16'hfe00;
			16'h81eb: y = 16'hfe00;
			16'h81ec: y = 16'hfe00;
			16'h81ed: y = 16'hfe00;
			16'h81ee: y = 16'hfe00;
			16'h81ef: y = 16'hfe00;
			16'h81f0: y = 16'hfe00;
			16'h81f1: y = 16'hfe00;
			16'h81f2: y = 16'hfe00;
			16'h81f3: y = 16'hfe00;
			16'h81f4: y = 16'hfe00;
			16'h81f5: y = 16'hfe00;
			16'h81f6: y = 16'hfe00;
			16'h81f7: y = 16'hfe00;
			16'h81f8: y = 16'hfe00;
			16'h81f9: y = 16'hfe00;
			16'h81fa: y = 16'hfe00;
			16'h81fb: y = 16'hfe00;
			16'h81fc: y = 16'hfe00;
			16'h81fd: y = 16'hfe00;
			16'h81fe: y = 16'hfe00;
			16'h81ff: y = 16'hfe00;
			16'h8200: y = 16'hfe00;
			16'h8201: y = 16'hfe00;
			16'h8202: y = 16'hfe00;
			16'h8203: y = 16'hfe00;
			16'h8204: y = 16'hfe00;
			16'h8205: y = 16'hfe00;
			16'h8206: y = 16'hfe00;
			16'h8207: y = 16'hfe00;
			16'h8208: y = 16'hfe00;
			16'h8209: y = 16'hfe00;
			16'h820a: y = 16'hfe00;
			16'h820b: y = 16'hfe00;
			16'h820c: y = 16'hfe00;
			16'h820d: y = 16'hfe00;
			16'h820e: y = 16'hfe00;
			16'h820f: y = 16'hfe00;
			16'h8210: y = 16'hfe00;
			16'h8211: y = 16'hfe00;
			16'h8212: y = 16'hfe00;
			16'h8213: y = 16'hfe00;
			16'h8214: y = 16'hfe00;
			16'h8215: y = 16'hfe00;
			16'h8216: y = 16'hfe00;
			16'h8217: y = 16'hfe00;
			16'h8218: y = 16'hfe00;
			16'h8219: y = 16'hfe00;
			16'h821a: y = 16'hfe00;
			16'h821b: y = 16'hfe00;
			16'h821c: y = 16'hfe00;
			16'h821d: y = 16'hfe00;
			16'h821e: y = 16'hfe00;
			16'h821f: y = 16'hfe00;
			16'h8220: y = 16'hfe00;
			16'h8221: y = 16'hfe00;
			16'h8222: y = 16'hfe00;
			16'h8223: y = 16'hfe00;
			16'h8224: y = 16'hfe00;
			16'h8225: y = 16'hfe00;
			16'h8226: y = 16'hfe00;
			16'h8227: y = 16'hfe00;
			16'h8228: y = 16'hfe00;
			16'h8229: y = 16'hfe00;
			16'h822a: y = 16'hfe00;
			16'h822b: y = 16'hfe00;
			16'h822c: y = 16'hfe00;
			16'h822d: y = 16'hfe00;
			16'h822e: y = 16'hfe00;
			16'h822f: y = 16'hfe00;
			16'h8230: y = 16'hfe00;
			16'h8231: y = 16'hfe00;
			16'h8232: y = 16'hfe00;
			16'h8233: y = 16'hfe00;
			16'h8234: y = 16'hfe00;
			16'h8235: y = 16'hfe00;
			16'h8236: y = 16'hfe00;
			16'h8237: y = 16'hfe00;
			16'h8238: y = 16'hfe00;
			16'h8239: y = 16'hfe00;
			16'h823a: y = 16'hfe00;
			16'h823b: y = 16'hfe00;
			16'h823c: y = 16'hfe00;
			16'h823d: y = 16'hfe00;
			16'h823e: y = 16'hfe00;
			16'h823f: y = 16'hfe00;
			16'h8240: y = 16'hfe00;
			16'h8241: y = 16'hfe00;
			16'h8242: y = 16'hfe00;
			16'h8243: y = 16'hfe00;
			16'h8244: y = 16'hfe00;
			16'h8245: y = 16'hfe00;
			16'h8246: y = 16'hfe00;
			16'h8247: y = 16'hfe00;
			16'h8248: y = 16'hfe00;
			16'h8249: y = 16'hfe00;
			16'h824a: y = 16'hfe00;
			16'h824b: y = 16'hfe00;
			16'h824c: y = 16'hfe00;
			16'h824d: y = 16'hfe00;
			16'h824e: y = 16'hfe00;
			16'h824f: y = 16'hfe00;
			16'h8250: y = 16'hfe00;
			16'h8251: y = 16'hfe00;
			16'h8252: y = 16'hfe00;
			16'h8253: y = 16'hfe00;
			16'h8254: y = 16'hfe00;
			16'h8255: y = 16'hfe00;
			16'h8256: y = 16'hfe00;
			16'h8257: y = 16'hfe00;
			16'h8258: y = 16'hfe00;
			16'h8259: y = 16'hfe00;
			16'h825a: y = 16'hfe00;
			16'h825b: y = 16'hfe00;
			16'h825c: y = 16'hfe00;
			16'h825d: y = 16'hfe00;
			16'h825e: y = 16'hfe00;
			16'h825f: y = 16'hfe00;
			16'h8260: y = 16'hfe00;
			16'h8261: y = 16'hfe00;
			16'h8262: y = 16'hfe00;
			16'h8263: y = 16'hfe00;
			16'h8264: y = 16'hfe00;
			16'h8265: y = 16'hfe00;
			16'h8266: y = 16'hfe00;
			16'h8267: y = 16'hfe00;
			16'h8268: y = 16'hfe00;
			16'h8269: y = 16'hfe00;
			16'h826a: y = 16'hfe00;
			16'h826b: y = 16'hfe00;
			16'h826c: y = 16'hfe00;
			16'h826d: y = 16'hfe00;
			16'h826e: y = 16'hfe00;
			16'h826f: y = 16'hfe00;
			16'h8270: y = 16'hfe00;
			16'h8271: y = 16'hfe00;
			16'h8272: y = 16'hfe00;
			16'h8273: y = 16'hfe00;
			16'h8274: y = 16'hfe00;
			16'h8275: y = 16'hfe00;
			16'h8276: y = 16'hfe00;
			16'h8277: y = 16'hfe00;
			16'h8278: y = 16'hfe00;
			16'h8279: y = 16'hfe00;
			16'h827a: y = 16'hfe00;
			16'h827b: y = 16'hfe00;
			16'h827c: y = 16'hfe00;
			16'h827d: y = 16'hfe00;
			16'h827e: y = 16'hfe00;
			16'h827f: y = 16'hfe00;
			16'h8280: y = 16'hfe00;
			16'h8281: y = 16'hfe00;
			16'h8282: y = 16'hfe00;
			16'h8283: y = 16'hfe00;
			16'h8284: y = 16'hfe00;
			16'h8285: y = 16'hfe00;
			16'h8286: y = 16'hfe00;
			16'h8287: y = 16'hfe00;
			16'h8288: y = 16'hfe00;
			16'h8289: y = 16'hfe00;
			16'h828a: y = 16'hfe00;
			16'h828b: y = 16'hfe00;
			16'h828c: y = 16'hfe00;
			16'h828d: y = 16'hfe00;
			16'h828e: y = 16'hfe00;
			16'h828f: y = 16'hfe00;
			16'h8290: y = 16'hfe00;
			16'h8291: y = 16'hfe00;
			16'h8292: y = 16'hfe00;
			16'h8293: y = 16'hfe00;
			16'h8294: y = 16'hfe00;
			16'h8295: y = 16'hfe00;
			16'h8296: y = 16'hfe00;
			16'h8297: y = 16'hfe00;
			16'h8298: y = 16'hfe00;
			16'h8299: y = 16'hfe00;
			16'h829a: y = 16'hfe00;
			16'h829b: y = 16'hfe00;
			16'h829c: y = 16'hfe00;
			16'h829d: y = 16'hfe00;
			16'h829e: y = 16'hfe00;
			16'h829f: y = 16'hfe00;
			16'h82a0: y = 16'hfe00;
			16'h82a1: y = 16'hfe00;
			16'h82a2: y = 16'hfe00;
			16'h82a3: y = 16'hfe00;
			16'h82a4: y = 16'hfe00;
			16'h82a5: y = 16'hfe00;
			16'h82a6: y = 16'hfe00;
			16'h82a7: y = 16'hfe00;
			16'h82a8: y = 16'hfe00;
			16'h82a9: y = 16'hfe00;
			16'h82aa: y = 16'hfe00;
			16'h82ab: y = 16'hfe00;
			16'h82ac: y = 16'hfe00;
			16'h82ad: y = 16'hfe00;
			16'h82ae: y = 16'hfe00;
			16'h82af: y = 16'hfe00;
			16'h82b0: y = 16'hfe00;
			16'h82b1: y = 16'hfe00;
			16'h82b2: y = 16'hfe00;
			16'h82b3: y = 16'hfe00;
			16'h82b4: y = 16'hfe00;
			16'h82b5: y = 16'hfe00;
			16'h82b6: y = 16'hfe00;
			16'h82b7: y = 16'hfe00;
			16'h82b8: y = 16'hfe00;
			16'h82b9: y = 16'hfe00;
			16'h82ba: y = 16'hfe00;
			16'h82bb: y = 16'hfe00;
			16'h82bc: y = 16'hfe00;
			16'h82bd: y = 16'hfe00;
			16'h82be: y = 16'hfe00;
			16'h82bf: y = 16'hfe00;
			16'h82c0: y = 16'hfe00;
			16'h82c1: y = 16'hfe00;
			16'h82c2: y = 16'hfe00;
			16'h82c3: y = 16'hfe00;
			16'h82c4: y = 16'hfe00;
			16'h82c5: y = 16'hfe00;
			16'h82c6: y = 16'hfe00;
			16'h82c7: y = 16'hfe00;
			16'h82c8: y = 16'hfe00;
			16'h82c9: y = 16'hfe00;
			16'h82ca: y = 16'hfe00;
			16'h82cb: y = 16'hfe00;
			16'h82cc: y = 16'hfe00;
			16'h82cd: y = 16'hfe00;
			16'h82ce: y = 16'hfe00;
			16'h82cf: y = 16'hfe00;
			16'h82d0: y = 16'hfe00;
			16'h82d1: y = 16'hfe00;
			16'h82d2: y = 16'hfe00;
			16'h82d3: y = 16'hfe00;
			16'h82d4: y = 16'hfe00;
			16'h82d5: y = 16'hfe00;
			16'h82d6: y = 16'hfe00;
			16'h82d7: y = 16'hfe00;
			16'h82d8: y = 16'hfe00;
			16'h82d9: y = 16'hfe00;
			16'h82da: y = 16'hfe00;
			16'h82db: y = 16'hfe00;
			16'h82dc: y = 16'hfe00;
			16'h82dd: y = 16'hfe00;
			16'h82de: y = 16'hfe00;
			16'h82df: y = 16'hfe00;
			16'h82e0: y = 16'hfe00;
			16'h82e1: y = 16'hfe00;
			16'h82e2: y = 16'hfe00;
			16'h82e3: y = 16'hfe00;
			16'h82e4: y = 16'hfe00;
			16'h82e5: y = 16'hfe00;
			16'h82e6: y = 16'hfe00;
			16'h82e7: y = 16'hfe00;
			16'h82e8: y = 16'hfe00;
			16'h82e9: y = 16'hfe00;
			16'h82ea: y = 16'hfe00;
			16'h82eb: y = 16'hfe00;
			16'h82ec: y = 16'hfe00;
			16'h82ed: y = 16'hfe00;
			16'h82ee: y = 16'hfe00;
			16'h82ef: y = 16'hfe00;
			16'h82f0: y = 16'hfe00;
			16'h82f1: y = 16'hfe00;
			16'h82f2: y = 16'hfe00;
			16'h82f3: y = 16'hfe00;
			16'h82f4: y = 16'hfe00;
			16'h82f5: y = 16'hfe00;
			16'h82f6: y = 16'hfe00;
			16'h82f7: y = 16'hfe00;
			16'h82f8: y = 16'hfe00;
			16'h82f9: y = 16'hfe00;
			16'h82fa: y = 16'hfe00;
			16'h82fb: y = 16'hfe00;
			16'h82fc: y = 16'hfe00;
			16'h82fd: y = 16'hfe00;
			16'h82fe: y = 16'hfe00;
			16'h82ff: y = 16'hfe00;
			16'h8300: y = 16'hfe00;
			16'h8301: y = 16'hfe00;
			16'h8302: y = 16'hfe00;
			16'h8303: y = 16'hfe00;
			16'h8304: y = 16'hfe00;
			16'h8305: y = 16'hfe00;
			16'h8306: y = 16'hfe00;
			16'h8307: y = 16'hfe00;
			16'h8308: y = 16'hfe00;
			16'h8309: y = 16'hfe00;
			16'h830a: y = 16'hfe00;
			16'h830b: y = 16'hfe00;
			16'h830c: y = 16'hfe00;
			16'h830d: y = 16'hfe00;
			16'h830e: y = 16'hfe00;
			16'h830f: y = 16'hfe00;
			16'h8310: y = 16'hfe00;
			16'h8311: y = 16'hfe00;
			16'h8312: y = 16'hfe00;
			16'h8313: y = 16'hfe00;
			16'h8314: y = 16'hfe00;
			16'h8315: y = 16'hfe00;
			16'h8316: y = 16'hfe00;
			16'h8317: y = 16'hfe00;
			16'h8318: y = 16'hfe00;
			16'h8319: y = 16'hfe00;
			16'h831a: y = 16'hfe00;
			16'h831b: y = 16'hfe00;
			16'h831c: y = 16'hfe00;
			16'h831d: y = 16'hfe00;
			16'h831e: y = 16'hfe00;
			16'h831f: y = 16'hfe00;
			16'h8320: y = 16'hfe00;
			16'h8321: y = 16'hfe00;
			16'h8322: y = 16'hfe00;
			16'h8323: y = 16'hfe00;
			16'h8324: y = 16'hfe00;
			16'h8325: y = 16'hfe00;
			16'h8326: y = 16'hfe00;
			16'h8327: y = 16'hfe00;
			16'h8328: y = 16'hfe00;
			16'h8329: y = 16'hfe00;
			16'h832a: y = 16'hfe00;
			16'h832b: y = 16'hfe00;
			16'h832c: y = 16'hfe00;
			16'h832d: y = 16'hfe00;
			16'h832e: y = 16'hfe00;
			16'h832f: y = 16'hfe00;
			16'h8330: y = 16'hfe00;
			16'h8331: y = 16'hfe00;
			16'h8332: y = 16'hfe00;
			16'h8333: y = 16'hfe00;
			16'h8334: y = 16'hfe00;
			16'h8335: y = 16'hfe00;
			16'h8336: y = 16'hfe00;
			16'h8337: y = 16'hfe00;
			16'h8338: y = 16'hfe00;
			16'h8339: y = 16'hfe00;
			16'h833a: y = 16'hfe00;
			16'h833b: y = 16'hfe00;
			16'h833c: y = 16'hfe00;
			16'h833d: y = 16'hfe00;
			16'h833e: y = 16'hfe00;
			16'h833f: y = 16'hfe00;
			16'h8340: y = 16'hfe00;
			16'h8341: y = 16'hfe00;
			16'h8342: y = 16'hfe00;
			16'h8343: y = 16'hfe00;
			16'h8344: y = 16'hfe00;
			16'h8345: y = 16'hfe00;
			16'h8346: y = 16'hfe00;
			16'h8347: y = 16'hfe00;
			16'h8348: y = 16'hfe00;
			16'h8349: y = 16'hfe00;
			16'h834a: y = 16'hfe00;
			16'h834b: y = 16'hfe00;
			16'h834c: y = 16'hfe00;
			16'h834d: y = 16'hfe00;
			16'h834e: y = 16'hfe00;
			16'h834f: y = 16'hfe00;
			16'h8350: y = 16'hfe00;
			16'h8351: y = 16'hfe00;
			16'h8352: y = 16'hfe00;
			16'h8353: y = 16'hfe00;
			16'h8354: y = 16'hfe00;
			16'h8355: y = 16'hfe00;
			16'h8356: y = 16'hfe00;
			16'h8357: y = 16'hfe00;
			16'h8358: y = 16'hfe00;
			16'h8359: y = 16'hfe00;
			16'h835a: y = 16'hfe00;
			16'h835b: y = 16'hfe00;
			16'h835c: y = 16'hfe00;
			16'h835d: y = 16'hfe00;
			16'h835e: y = 16'hfe00;
			16'h835f: y = 16'hfe00;
			16'h8360: y = 16'hfe00;
			16'h8361: y = 16'hfe00;
			16'h8362: y = 16'hfe00;
			16'h8363: y = 16'hfe00;
			16'h8364: y = 16'hfe00;
			16'h8365: y = 16'hfe00;
			16'h8366: y = 16'hfe00;
			16'h8367: y = 16'hfe00;
			16'h8368: y = 16'hfe00;
			16'h8369: y = 16'hfe00;
			16'h836a: y = 16'hfe00;
			16'h836b: y = 16'hfe00;
			16'h836c: y = 16'hfe00;
			16'h836d: y = 16'hfe00;
			16'h836e: y = 16'hfe00;
			16'h836f: y = 16'hfe00;
			16'h8370: y = 16'hfe00;
			16'h8371: y = 16'hfe00;
			16'h8372: y = 16'hfe00;
			16'h8373: y = 16'hfe00;
			16'h8374: y = 16'hfe00;
			16'h8375: y = 16'hfe00;
			16'h8376: y = 16'hfe00;
			16'h8377: y = 16'hfe00;
			16'h8378: y = 16'hfe00;
			16'h8379: y = 16'hfe00;
			16'h837a: y = 16'hfe00;
			16'h837b: y = 16'hfe00;
			16'h837c: y = 16'hfe00;
			16'h837d: y = 16'hfe00;
			16'h837e: y = 16'hfe00;
			16'h837f: y = 16'hfe00;
			16'h8380: y = 16'hfe00;
			16'h8381: y = 16'hfe00;
			16'h8382: y = 16'hfe00;
			16'h8383: y = 16'hfe00;
			16'h8384: y = 16'hfe00;
			16'h8385: y = 16'hfe00;
			16'h8386: y = 16'hfe00;
			16'h8387: y = 16'hfe00;
			16'h8388: y = 16'hfe00;
			16'h8389: y = 16'hfe00;
			16'h838a: y = 16'hfe00;
			16'h838b: y = 16'hfe00;
			16'h838c: y = 16'hfe00;
			16'h838d: y = 16'hfe00;
			16'h838e: y = 16'hfe00;
			16'h838f: y = 16'hfe00;
			16'h8390: y = 16'hfe00;
			16'h8391: y = 16'hfe00;
			16'h8392: y = 16'hfe00;
			16'h8393: y = 16'hfe00;
			16'h8394: y = 16'hfe00;
			16'h8395: y = 16'hfe00;
			16'h8396: y = 16'hfe00;
			16'h8397: y = 16'hfe00;
			16'h8398: y = 16'hfe00;
			16'h8399: y = 16'hfe00;
			16'h839a: y = 16'hfe00;
			16'h839b: y = 16'hfe00;
			16'h839c: y = 16'hfe00;
			16'h839d: y = 16'hfe00;
			16'h839e: y = 16'hfe00;
			16'h839f: y = 16'hfe00;
			16'h83a0: y = 16'hfe00;
			16'h83a1: y = 16'hfe00;
			16'h83a2: y = 16'hfe00;
			16'h83a3: y = 16'hfe00;
			16'h83a4: y = 16'hfe00;
			16'h83a5: y = 16'hfe00;
			16'h83a6: y = 16'hfe00;
			16'h83a7: y = 16'hfe00;
			16'h83a8: y = 16'hfe00;
			16'h83a9: y = 16'hfe00;
			16'h83aa: y = 16'hfe00;
			16'h83ab: y = 16'hfe00;
			16'h83ac: y = 16'hfe00;
			16'h83ad: y = 16'hfe00;
			16'h83ae: y = 16'hfe00;
			16'h83af: y = 16'hfe00;
			16'h83b0: y = 16'hfe00;
			16'h83b1: y = 16'hfe00;
			16'h83b2: y = 16'hfe00;
			16'h83b3: y = 16'hfe00;
			16'h83b4: y = 16'hfe00;
			16'h83b5: y = 16'hfe00;
			16'h83b6: y = 16'hfe00;
			16'h83b7: y = 16'hfe00;
			16'h83b8: y = 16'hfe00;
			16'h83b9: y = 16'hfe00;
			16'h83ba: y = 16'hfe00;
			16'h83bb: y = 16'hfe00;
			16'h83bc: y = 16'hfe00;
			16'h83bd: y = 16'hfe00;
			16'h83be: y = 16'hfe00;
			16'h83bf: y = 16'hfe00;
			16'h83c0: y = 16'hfe00;
			16'h83c1: y = 16'hfe00;
			16'h83c2: y = 16'hfe00;
			16'h83c3: y = 16'hfe00;
			16'h83c4: y = 16'hfe00;
			16'h83c5: y = 16'hfe00;
			16'h83c6: y = 16'hfe00;
			16'h83c7: y = 16'hfe00;
			16'h83c8: y = 16'hfe00;
			16'h83c9: y = 16'hfe00;
			16'h83ca: y = 16'hfe00;
			16'h83cb: y = 16'hfe00;
			16'h83cc: y = 16'hfe00;
			16'h83cd: y = 16'hfe00;
			16'h83ce: y = 16'hfe00;
			16'h83cf: y = 16'hfe00;
			16'h83d0: y = 16'hfe00;
			16'h83d1: y = 16'hfe00;
			16'h83d2: y = 16'hfe00;
			16'h83d3: y = 16'hfe00;
			16'h83d4: y = 16'hfe00;
			16'h83d5: y = 16'hfe00;
			16'h83d6: y = 16'hfe00;
			16'h83d7: y = 16'hfe00;
			16'h83d8: y = 16'hfe00;
			16'h83d9: y = 16'hfe00;
			16'h83da: y = 16'hfe00;
			16'h83db: y = 16'hfe00;
			16'h83dc: y = 16'hfe00;
			16'h83dd: y = 16'hfe00;
			16'h83de: y = 16'hfe00;
			16'h83df: y = 16'hfe00;
			16'h83e0: y = 16'hfe00;
			16'h83e1: y = 16'hfe00;
			16'h83e2: y = 16'hfe00;
			16'h83e3: y = 16'hfe00;
			16'h83e4: y = 16'hfe00;
			16'h83e5: y = 16'hfe00;
			16'h83e6: y = 16'hfe00;
			16'h83e7: y = 16'hfe00;
			16'h83e8: y = 16'hfe00;
			16'h83e9: y = 16'hfe00;
			16'h83ea: y = 16'hfe00;
			16'h83eb: y = 16'hfe00;
			16'h83ec: y = 16'hfe00;
			16'h83ed: y = 16'hfe00;
			16'h83ee: y = 16'hfe00;
			16'h83ef: y = 16'hfe00;
			16'h83f0: y = 16'hfe00;
			16'h83f1: y = 16'hfe00;
			16'h83f2: y = 16'hfe00;
			16'h83f3: y = 16'hfe00;
			16'h83f4: y = 16'hfe00;
			16'h83f5: y = 16'hfe00;
			16'h83f6: y = 16'hfe00;
			16'h83f7: y = 16'hfe00;
			16'h83f8: y = 16'hfe00;
			16'h83f9: y = 16'hfe00;
			16'h83fa: y = 16'hfe00;
			16'h83fb: y = 16'hfe00;
			16'h83fc: y = 16'hfe00;
			16'h83fd: y = 16'hfe00;
			16'h83fe: y = 16'hfe00;
			16'h83ff: y = 16'hfe00;
			16'h8400: y = 16'hfe00;
			16'h8401: y = 16'hfe00;
			16'h8402: y = 16'hfe00;
			16'h8403: y = 16'hfe00;
			16'h8404: y = 16'hfe00;
			16'h8405: y = 16'hfe00;
			16'h8406: y = 16'hfe00;
			16'h8407: y = 16'hfe00;
			16'h8408: y = 16'hfe00;
			16'h8409: y = 16'hfe00;
			16'h840a: y = 16'hfe00;
			16'h840b: y = 16'hfe00;
			16'h840c: y = 16'hfe00;
			16'h840d: y = 16'hfe00;
			16'h840e: y = 16'hfe00;
			16'h840f: y = 16'hfe00;
			16'h8410: y = 16'hfe00;
			16'h8411: y = 16'hfe00;
			16'h8412: y = 16'hfe00;
			16'h8413: y = 16'hfe00;
			16'h8414: y = 16'hfe00;
			16'h8415: y = 16'hfe00;
			16'h8416: y = 16'hfe00;
			16'h8417: y = 16'hfe00;
			16'h8418: y = 16'hfe00;
			16'h8419: y = 16'hfe00;
			16'h841a: y = 16'hfe00;
			16'h841b: y = 16'hfe00;
			16'h841c: y = 16'hfe00;
			16'h841d: y = 16'hfe00;
			16'h841e: y = 16'hfe00;
			16'h841f: y = 16'hfe00;
			16'h8420: y = 16'hfe00;
			16'h8421: y = 16'hfe00;
			16'h8422: y = 16'hfe00;
			16'h8423: y = 16'hfe00;
			16'h8424: y = 16'hfe00;
			16'h8425: y = 16'hfe00;
			16'h8426: y = 16'hfe00;
			16'h8427: y = 16'hfe00;
			16'h8428: y = 16'hfe00;
			16'h8429: y = 16'hfe00;
			16'h842a: y = 16'hfe00;
			16'h842b: y = 16'hfe00;
			16'h842c: y = 16'hfe00;
			16'h842d: y = 16'hfe00;
			16'h842e: y = 16'hfe00;
			16'h842f: y = 16'hfe00;
			16'h8430: y = 16'hfe00;
			16'h8431: y = 16'hfe00;
			16'h8432: y = 16'hfe00;
			16'h8433: y = 16'hfe00;
			16'h8434: y = 16'hfe00;
			16'h8435: y = 16'hfe00;
			16'h8436: y = 16'hfe00;
			16'h8437: y = 16'hfe00;
			16'h8438: y = 16'hfe00;
			16'h8439: y = 16'hfe00;
			16'h843a: y = 16'hfe00;
			16'h843b: y = 16'hfe00;
			16'h843c: y = 16'hfe00;
			16'h843d: y = 16'hfe00;
			16'h843e: y = 16'hfe00;
			16'h843f: y = 16'hfe00;
			16'h8440: y = 16'hfe00;
			16'h8441: y = 16'hfe00;
			16'h8442: y = 16'hfe00;
			16'h8443: y = 16'hfe00;
			16'h8444: y = 16'hfe00;
			16'h8445: y = 16'hfe00;
			16'h8446: y = 16'hfe00;
			16'h8447: y = 16'hfe00;
			16'h8448: y = 16'hfe00;
			16'h8449: y = 16'hfe00;
			16'h844a: y = 16'hfe00;
			16'h844b: y = 16'hfe00;
			16'h844c: y = 16'hfe00;
			16'h844d: y = 16'hfe00;
			16'h844e: y = 16'hfe00;
			16'h844f: y = 16'hfe00;
			16'h8450: y = 16'hfe00;
			16'h8451: y = 16'hfe00;
			16'h8452: y = 16'hfe00;
			16'h8453: y = 16'hfe00;
			16'h8454: y = 16'hfe00;
			16'h8455: y = 16'hfe00;
			16'h8456: y = 16'hfe00;
			16'h8457: y = 16'hfe00;
			16'h8458: y = 16'hfe00;
			16'h8459: y = 16'hfe00;
			16'h845a: y = 16'hfe00;
			16'h845b: y = 16'hfe00;
			16'h845c: y = 16'hfe00;
			16'h845d: y = 16'hfe00;
			16'h845e: y = 16'hfe00;
			16'h845f: y = 16'hfe00;
			16'h8460: y = 16'hfe00;
			16'h8461: y = 16'hfe00;
			16'h8462: y = 16'hfe00;
			16'h8463: y = 16'hfe00;
			16'h8464: y = 16'hfe00;
			16'h8465: y = 16'hfe00;
			16'h8466: y = 16'hfe00;
			16'h8467: y = 16'hfe00;
			16'h8468: y = 16'hfe00;
			16'h8469: y = 16'hfe00;
			16'h846a: y = 16'hfe00;
			16'h846b: y = 16'hfe00;
			16'h846c: y = 16'hfe00;
			16'h846d: y = 16'hfe00;
			16'h846e: y = 16'hfe00;
			16'h846f: y = 16'hfe00;
			16'h8470: y = 16'hfe00;
			16'h8471: y = 16'hfe00;
			16'h8472: y = 16'hfe00;
			16'h8473: y = 16'hfe00;
			16'h8474: y = 16'hfe00;
			16'h8475: y = 16'hfe00;
			16'h8476: y = 16'hfe00;
			16'h8477: y = 16'hfe00;
			16'h8478: y = 16'hfe00;
			16'h8479: y = 16'hfe00;
			16'h847a: y = 16'hfe00;
			16'h847b: y = 16'hfe00;
			16'h847c: y = 16'hfe00;
			16'h847d: y = 16'hfe00;
			16'h847e: y = 16'hfe00;
			16'h847f: y = 16'hfe00;
			16'h8480: y = 16'hfe00;
			16'h8481: y = 16'hfe00;
			16'h8482: y = 16'hfe00;
			16'h8483: y = 16'hfe00;
			16'h8484: y = 16'hfe00;
			16'h8485: y = 16'hfe00;
			16'h8486: y = 16'hfe00;
			16'h8487: y = 16'hfe00;
			16'h8488: y = 16'hfe00;
			16'h8489: y = 16'hfe00;
			16'h848a: y = 16'hfe00;
			16'h848b: y = 16'hfe00;
			16'h848c: y = 16'hfe00;
			16'h848d: y = 16'hfe00;
			16'h848e: y = 16'hfe00;
			16'h848f: y = 16'hfe00;
			16'h8490: y = 16'hfe00;
			16'h8491: y = 16'hfe00;
			16'h8492: y = 16'hfe00;
			16'h8493: y = 16'hfe00;
			16'h8494: y = 16'hfe00;
			16'h8495: y = 16'hfe00;
			16'h8496: y = 16'hfe00;
			16'h8497: y = 16'hfe00;
			16'h8498: y = 16'hfe00;
			16'h8499: y = 16'hfe00;
			16'h849a: y = 16'hfe00;
			16'h849b: y = 16'hfe00;
			16'h849c: y = 16'hfe00;
			16'h849d: y = 16'hfe00;
			16'h849e: y = 16'hfe00;
			16'h849f: y = 16'hfe00;
			16'h84a0: y = 16'hfe00;
			16'h84a1: y = 16'hfe00;
			16'h84a2: y = 16'hfe00;
			16'h84a3: y = 16'hfe00;
			16'h84a4: y = 16'hfe00;
			16'h84a5: y = 16'hfe00;
			16'h84a6: y = 16'hfe00;
			16'h84a7: y = 16'hfe00;
			16'h84a8: y = 16'hfe00;
			16'h84a9: y = 16'hfe00;
			16'h84aa: y = 16'hfe00;
			16'h84ab: y = 16'hfe00;
			16'h84ac: y = 16'hfe00;
			16'h84ad: y = 16'hfe00;
			16'h84ae: y = 16'hfe00;
			16'h84af: y = 16'hfe00;
			16'h84b0: y = 16'hfe00;
			16'h84b1: y = 16'hfe00;
			16'h84b2: y = 16'hfe00;
			16'h84b3: y = 16'hfe00;
			16'h84b4: y = 16'hfe00;
			16'h84b5: y = 16'hfe00;
			16'h84b6: y = 16'hfe00;
			16'h84b7: y = 16'hfe00;
			16'h84b8: y = 16'hfe00;
			16'h84b9: y = 16'hfe00;
			16'h84ba: y = 16'hfe00;
			16'h84bb: y = 16'hfe00;
			16'h84bc: y = 16'hfe00;
			16'h84bd: y = 16'hfe00;
			16'h84be: y = 16'hfe00;
			16'h84bf: y = 16'hfe00;
			16'h84c0: y = 16'hfe00;
			16'h84c1: y = 16'hfe00;
			16'h84c2: y = 16'hfe00;
			16'h84c3: y = 16'hfe00;
			16'h84c4: y = 16'hfe00;
			16'h84c5: y = 16'hfe00;
			16'h84c6: y = 16'hfe00;
			16'h84c7: y = 16'hfe00;
			16'h84c8: y = 16'hfe00;
			16'h84c9: y = 16'hfe00;
			16'h84ca: y = 16'hfe00;
			16'h84cb: y = 16'hfe00;
			16'h84cc: y = 16'hfe00;
			16'h84cd: y = 16'hfe00;
			16'h84ce: y = 16'hfe00;
			16'h84cf: y = 16'hfe00;
			16'h84d0: y = 16'hfe00;
			16'h84d1: y = 16'hfe00;
			16'h84d2: y = 16'hfe00;
			16'h84d3: y = 16'hfe00;
			16'h84d4: y = 16'hfe00;
			16'h84d5: y = 16'hfe00;
			16'h84d6: y = 16'hfe00;
			16'h84d7: y = 16'hfe00;
			16'h84d8: y = 16'hfe00;
			16'h84d9: y = 16'hfe00;
			16'h84da: y = 16'hfe00;
			16'h84db: y = 16'hfe00;
			16'h84dc: y = 16'hfe00;
			16'h84dd: y = 16'hfe00;
			16'h84de: y = 16'hfe00;
			16'h84df: y = 16'hfe00;
			16'h84e0: y = 16'hfe00;
			16'h84e1: y = 16'hfe00;
			16'h84e2: y = 16'hfe00;
			16'h84e3: y = 16'hfe00;
			16'h84e4: y = 16'hfe00;
			16'h84e5: y = 16'hfe00;
			16'h84e6: y = 16'hfe00;
			16'h84e7: y = 16'hfe00;
			16'h84e8: y = 16'hfe00;
			16'h84e9: y = 16'hfe00;
			16'h84ea: y = 16'hfe00;
			16'h84eb: y = 16'hfe00;
			16'h84ec: y = 16'hfe00;
			16'h84ed: y = 16'hfe00;
			16'h84ee: y = 16'hfe00;
			16'h84ef: y = 16'hfe00;
			16'h84f0: y = 16'hfe00;
			16'h84f1: y = 16'hfe00;
			16'h84f2: y = 16'hfe00;
			16'h84f3: y = 16'hfe00;
			16'h84f4: y = 16'hfe00;
			16'h84f5: y = 16'hfe00;
			16'h84f6: y = 16'hfe00;
			16'h84f7: y = 16'hfe00;
			16'h84f8: y = 16'hfe00;
			16'h84f9: y = 16'hfe00;
			16'h84fa: y = 16'hfe00;
			16'h84fb: y = 16'hfe00;
			16'h84fc: y = 16'hfe00;
			16'h84fd: y = 16'hfe00;
			16'h84fe: y = 16'hfe00;
			16'h84ff: y = 16'hfe00;
			16'h8500: y = 16'hfe00;
			16'h8501: y = 16'hfe00;
			16'h8502: y = 16'hfe00;
			16'h8503: y = 16'hfe00;
			16'h8504: y = 16'hfe00;
			16'h8505: y = 16'hfe00;
			16'h8506: y = 16'hfe00;
			16'h8507: y = 16'hfe00;
			16'h8508: y = 16'hfe00;
			16'h8509: y = 16'hfe00;
			16'h850a: y = 16'hfe00;
			16'h850b: y = 16'hfe00;
			16'h850c: y = 16'hfe00;
			16'h850d: y = 16'hfe00;
			16'h850e: y = 16'hfe00;
			16'h850f: y = 16'hfe00;
			16'h8510: y = 16'hfe00;
			16'h8511: y = 16'hfe00;
			16'h8512: y = 16'hfe00;
			16'h8513: y = 16'hfe00;
			16'h8514: y = 16'hfe00;
			16'h8515: y = 16'hfe00;
			16'h8516: y = 16'hfe00;
			16'h8517: y = 16'hfe00;
			16'h8518: y = 16'hfe00;
			16'h8519: y = 16'hfe00;
			16'h851a: y = 16'hfe00;
			16'h851b: y = 16'hfe00;
			16'h851c: y = 16'hfe00;
			16'h851d: y = 16'hfe00;
			16'h851e: y = 16'hfe00;
			16'h851f: y = 16'hfe00;
			16'h8520: y = 16'hfe00;
			16'h8521: y = 16'hfe00;
			16'h8522: y = 16'hfe00;
			16'h8523: y = 16'hfe00;
			16'h8524: y = 16'hfe00;
			16'h8525: y = 16'hfe00;
			16'h8526: y = 16'hfe00;
			16'h8527: y = 16'hfe00;
			16'h8528: y = 16'hfe00;
			16'h8529: y = 16'hfe00;
			16'h852a: y = 16'hfe00;
			16'h852b: y = 16'hfe00;
			16'h852c: y = 16'hfe00;
			16'h852d: y = 16'hfe00;
			16'h852e: y = 16'hfe00;
			16'h852f: y = 16'hfe00;
			16'h8530: y = 16'hfe00;
			16'h8531: y = 16'hfe00;
			16'h8532: y = 16'hfe00;
			16'h8533: y = 16'hfe00;
			16'h8534: y = 16'hfe00;
			16'h8535: y = 16'hfe00;
			16'h8536: y = 16'hfe00;
			16'h8537: y = 16'hfe00;
			16'h8538: y = 16'hfe00;
			16'h8539: y = 16'hfe00;
			16'h853a: y = 16'hfe00;
			16'h853b: y = 16'hfe00;
			16'h853c: y = 16'hfe00;
			16'h853d: y = 16'hfe00;
			16'h853e: y = 16'hfe00;
			16'h853f: y = 16'hfe00;
			16'h8540: y = 16'hfe00;
			16'h8541: y = 16'hfe00;
			16'h8542: y = 16'hfe00;
			16'h8543: y = 16'hfe00;
			16'h8544: y = 16'hfe00;
			16'h8545: y = 16'hfe00;
			16'h8546: y = 16'hfe00;
			16'h8547: y = 16'hfe00;
			16'h8548: y = 16'hfe00;
			16'h8549: y = 16'hfe00;
			16'h854a: y = 16'hfe00;
			16'h854b: y = 16'hfe00;
			16'h854c: y = 16'hfe00;
			16'h854d: y = 16'hfe00;
			16'h854e: y = 16'hfe00;
			16'h854f: y = 16'hfe00;
			16'h8550: y = 16'hfe00;
			16'h8551: y = 16'hfe00;
			16'h8552: y = 16'hfe00;
			16'h8553: y = 16'hfe00;
			16'h8554: y = 16'hfe00;
			16'h8555: y = 16'hfe00;
			16'h8556: y = 16'hfe00;
			16'h8557: y = 16'hfe00;
			16'h8558: y = 16'hfe00;
			16'h8559: y = 16'hfe00;
			16'h855a: y = 16'hfe00;
			16'h855b: y = 16'hfe00;
			16'h855c: y = 16'hfe00;
			16'h855d: y = 16'hfe00;
			16'h855e: y = 16'hfe00;
			16'h855f: y = 16'hfe00;
			16'h8560: y = 16'hfe00;
			16'h8561: y = 16'hfe00;
			16'h8562: y = 16'hfe00;
			16'h8563: y = 16'hfe00;
			16'h8564: y = 16'hfe00;
			16'h8565: y = 16'hfe00;
			16'h8566: y = 16'hfe00;
			16'h8567: y = 16'hfe00;
			16'h8568: y = 16'hfe00;
			16'h8569: y = 16'hfe00;
			16'h856a: y = 16'hfe00;
			16'h856b: y = 16'hfe00;
			16'h856c: y = 16'hfe00;
			16'h856d: y = 16'hfe00;
			16'h856e: y = 16'hfe00;
			16'h856f: y = 16'hfe00;
			16'h8570: y = 16'hfe00;
			16'h8571: y = 16'hfe00;
			16'h8572: y = 16'hfe00;
			16'h8573: y = 16'hfe00;
			16'h8574: y = 16'hfe00;
			16'h8575: y = 16'hfe00;
			16'h8576: y = 16'hfe00;
			16'h8577: y = 16'hfe00;
			16'h8578: y = 16'hfe00;
			16'h8579: y = 16'hfe00;
			16'h857a: y = 16'hfe00;
			16'h857b: y = 16'hfe00;
			16'h857c: y = 16'hfe00;
			16'h857d: y = 16'hfe00;
			16'h857e: y = 16'hfe00;
			16'h857f: y = 16'hfe00;
			16'h8580: y = 16'hfe00;
			16'h8581: y = 16'hfe00;
			16'h8582: y = 16'hfe00;
			16'h8583: y = 16'hfe00;
			16'h8584: y = 16'hfe00;
			16'h8585: y = 16'hfe00;
			16'h8586: y = 16'hfe00;
			16'h8587: y = 16'hfe00;
			16'h8588: y = 16'hfe00;
			16'h8589: y = 16'hfe00;
			16'h858a: y = 16'hfe00;
			16'h858b: y = 16'hfe00;
			16'h858c: y = 16'hfe00;
			16'h858d: y = 16'hfe00;
			16'h858e: y = 16'hfe00;
			16'h858f: y = 16'hfe00;
			16'h8590: y = 16'hfe00;
			16'h8591: y = 16'hfe00;
			16'h8592: y = 16'hfe00;
			16'h8593: y = 16'hfe00;
			16'h8594: y = 16'hfe00;
			16'h8595: y = 16'hfe00;
			16'h8596: y = 16'hfe00;
			16'h8597: y = 16'hfe00;
			16'h8598: y = 16'hfe00;
			16'h8599: y = 16'hfe00;
			16'h859a: y = 16'hfe00;
			16'h859b: y = 16'hfe00;
			16'h859c: y = 16'hfe00;
			16'h859d: y = 16'hfe00;
			16'h859e: y = 16'hfe00;
			16'h859f: y = 16'hfe00;
			16'h85a0: y = 16'hfe00;
			16'h85a1: y = 16'hfe00;
			16'h85a2: y = 16'hfe00;
			16'h85a3: y = 16'hfe00;
			16'h85a4: y = 16'hfe00;
			16'h85a5: y = 16'hfe00;
			16'h85a6: y = 16'hfe00;
			16'h85a7: y = 16'hfe00;
			16'h85a8: y = 16'hfe00;
			16'h85a9: y = 16'hfe00;
			16'h85aa: y = 16'hfe00;
			16'h85ab: y = 16'hfe00;
			16'h85ac: y = 16'hfe00;
			16'h85ad: y = 16'hfe00;
			16'h85ae: y = 16'hfe00;
			16'h85af: y = 16'hfe00;
			16'h85b0: y = 16'hfe00;
			16'h85b1: y = 16'hfe00;
			16'h85b2: y = 16'hfe00;
			16'h85b3: y = 16'hfe00;
			16'h85b4: y = 16'hfe00;
			16'h85b5: y = 16'hfe00;
			16'h85b6: y = 16'hfe00;
			16'h85b7: y = 16'hfe00;
			16'h85b8: y = 16'hfe00;
			16'h85b9: y = 16'hfe00;
			16'h85ba: y = 16'hfe00;
			16'h85bb: y = 16'hfe00;
			16'h85bc: y = 16'hfe00;
			16'h85bd: y = 16'hfe00;
			16'h85be: y = 16'hfe00;
			16'h85bf: y = 16'hfe00;
			16'h85c0: y = 16'hfe00;
			16'h85c1: y = 16'hfe00;
			16'h85c2: y = 16'hfe00;
			16'h85c3: y = 16'hfe00;
			16'h85c4: y = 16'hfe00;
			16'h85c5: y = 16'hfe00;
			16'h85c6: y = 16'hfe00;
			16'h85c7: y = 16'hfe00;
			16'h85c8: y = 16'hfe00;
			16'h85c9: y = 16'hfe00;
			16'h85ca: y = 16'hfe00;
			16'h85cb: y = 16'hfe00;
			16'h85cc: y = 16'hfe00;
			16'h85cd: y = 16'hfe00;
			16'h85ce: y = 16'hfe00;
			16'h85cf: y = 16'hfe00;
			16'h85d0: y = 16'hfe00;
			16'h85d1: y = 16'hfe00;
			16'h85d2: y = 16'hfe00;
			16'h85d3: y = 16'hfe00;
			16'h85d4: y = 16'hfe00;
			16'h85d5: y = 16'hfe00;
			16'h85d6: y = 16'hfe00;
			16'h85d7: y = 16'hfe00;
			16'h85d8: y = 16'hfe00;
			16'h85d9: y = 16'hfe00;
			16'h85da: y = 16'hfe00;
			16'h85db: y = 16'hfe00;
			16'h85dc: y = 16'hfe00;
			16'h85dd: y = 16'hfe00;
			16'h85de: y = 16'hfe00;
			16'h85df: y = 16'hfe00;
			16'h85e0: y = 16'hfe00;
			16'h85e1: y = 16'hfe00;
			16'h85e2: y = 16'hfe00;
			16'h85e3: y = 16'hfe00;
			16'h85e4: y = 16'hfe00;
			16'h85e5: y = 16'hfe00;
			16'h85e6: y = 16'hfe00;
			16'h85e7: y = 16'hfe00;
			16'h85e8: y = 16'hfe00;
			16'h85e9: y = 16'hfe00;
			16'h85ea: y = 16'hfe00;
			16'h85eb: y = 16'hfe00;
			16'h85ec: y = 16'hfe00;
			16'h85ed: y = 16'hfe00;
			16'h85ee: y = 16'hfe00;
			16'h85ef: y = 16'hfe00;
			16'h85f0: y = 16'hfe00;
			16'h85f1: y = 16'hfe00;
			16'h85f2: y = 16'hfe00;
			16'h85f3: y = 16'hfe00;
			16'h85f4: y = 16'hfe00;
			16'h85f5: y = 16'hfe00;
			16'h85f6: y = 16'hfe00;
			16'h85f7: y = 16'hfe00;
			16'h85f8: y = 16'hfe00;
			16'h85f9: y = 16'hfe00;
			16'h85fa: y = 16'hfe00;
			16'h85fb: y = 16'hfe00;
			16'h85fc: y = 16'hfe00;
			16'h85fd: y = 16'hfe00;
			16'h85fe: y = 16'hfe00;
			16'h85ff: y = 16'hfe00;
			16'h8600: y = 16'hfe00;
			16'h8601: y = 16'hfe00;
			16'h8602: y = 16'hfe00;
			16'h8603: y = 16'hfe00;
			16'h8604: y = 16'hfe00;
			16'h8605: y = 16'hfe00;
			16'h8606: y = 16'hfe00;
			16'h8607: y = 16'hfe00;
			16'h8608: y = 16'hfe00;
			16'h8609: y = 16'hfe00;
			16'h860a: y = 16'hfe00;
			16'h860b: y = 16'hfe00;
			16'h860c: y = 16'hfe00;
			16'h860d: y = 16'hfe00;
			16'h860e: y = 16'hfe00;
			16'h860f: y = 16'hfe00;
			16'h8610: y = 16'hfe00;
			16'h8611: y = 16'hfe00;
			16'h8612: y = 16'hfe00;
			16'h8613: y = 16'hfe00;
			16'h8614: y = 16'hfe00;
			16'h8615: y = 16'hfe00;
			16'h8616: y = 16'hfe00;
			16'h8617: y = 16'hfe00;
			16'h8618: y = 16'hfe00;
			16'h8619: y = 16'hfe00;
			16'h861a: y = 16'hfe00;
			16'h861b: y = 16'hfe00;
			16'h861c: y = 16'hfe00;
			16'h861d: y = 16'hfe00;
			16'h861e: y = 16'hfe00;
			16'h861f: y = 16'hfe00;
			16'h8620: y = 16'hfe00;
			16'h8621: y = 16'hfe00;
			16'h8622: y = 16'hfe00;
			16'h8623: y = 16'hfe00;
			16'h8624: y = 16'hfe00;
			16'h8625: y = 16'hfe00;
			16'h8626: y = 16'hfe00;
			16'h8627: y = 16'hfe00;
			16'h8628: y = 16'hfe00;
			16'h8629: y = 16'hfe00;
			16'h862a: y = 16'hfe00;
			16'h862b: y = 16'hfe00;
			16'h862c: y = 16'hfe00;
			16'h862d: y = 16'hfe00;
			16'h862e: y = 16'hfe00;
			16'h862f: y = 16'hfe00;
			16'h8630: y = 16'hfe00;
			16'h8631: y = 16'hfe00;
			16'h8632: y = 16'hfe00;
			16'h8633: y = 16'hfe00;
			16'h8634: y = 16'hfe00;
			16'h8635: y = 16'hfe00;
			16'h8636: y = 16'hfe00;
			16'h8637: y = 16'hfe00;
			16'h8638: y = 16'hfe00;
			16'h8639: y = 16'hfe00;
			16'h863a: y = 16'hfe00;
			16'h863b: y = 16'hfe00;
			16'h863c: y = 16'hfe00;
			16'h863d: y = 16'hfe00;
			16'h863e: y = 16'hfe00;
			16'h863f: y = 16'hfe00;
			16'h8640: y = 16'hfe00;
			16'h8641: y = 16'hfe00;
			16'h8642: y = 16'hfe00;
			16'h8643: y = 16'hfe00;
			16'h8644: y = 16'hfe00;
			16'h8645: y = 16'hfe00;
			16'h8646: y = 16'hfe00;
			16'h8647: y = 16'hfe00;
			16'h8648: y = 16'hfe00;
			16'h8649: y = 16'hfe00;
			16'h864a: y = 16'hfe00;
			16'h864b: y = 16'hfe00;
			16'h864c: y = 16'hfe00;
			16'h864d: y = 16'hfe00;
			16'h864e: y = 16'hfe00;
			16'h864f: y = 16'hfe00;
			16'h8650: y = 16'hfe00;
			16'h8651: y = 16'hfe00;
			16'h8652: y = 16'hfe00;
			16'h8653: y = 16'hfe00;
			16'h8654: y = 16'hfe00;
			16'h8655: y = 16'hfe00;
			16'h8656: y = 16'hfe00;
			16'h8657: y = 16'hfe00;
			16'h8658: y = 16'hfe00;
			16'h8659: y = 16'hfe00;
			16'h865a: y = 16'hfe00;
			16'h865b: y = 16'hfe00;
			16'h865c: y = 16'hfe00;
			16'h865d: y = 16'hfe00;
			16'h865e: y = 16'hfe00;
			16'h865f: y = 16'hfe00;
			16'h8660: y = 16'hfe00;
			16'h8661: y = 16'hfe00;
			16'h8662: y = 16'hfe00;
			16'h8663: y = 16'hfe00;
			16'h8664: y = 16'hfe00;
			16'h8665: y = 16'hfe00;
			16'h8666: y = 16'hfe00;
			16'h8667: y = 16'hfe00;
			16'h8668: y = 16'hfe00;
			16'h8669: y = 16'hfe00;
			16'h866a: y = 16'hfe00;
			16'h866b: y = 16'hfe00;
			16'h866c: y = 16'hfe00;
			16'h866d: y = 16'hfe00;
			16'h866e: y = 16'hfe00;
			16'h866f: y = 16'hfe00;
			16'h8670: y = 16'hfe00;
			16'h8671: y = 16'hfe00;
			16'h8672: y = 16'hfe00;
			16'h8673: y = 16'hfe00;
			16'h8674: y = 16'hfe00;
			16'h8675: y = 16'hfe00;
			16'h8676: y = 16'hfe00;
			16'h8677: y = 16'hfe00;
			16'h8678: y = 16'hfe00;
			16'h8679: y = 16'hfe00;
			16'h867a: y = 16'hfe00;
			16'h867b: y = 16'hfe00;
			16'h867c: y = 16'hfe00;
			16'h867d: y = 16'hfe00;
			16'h867e: y = 16'hfe00;
			16'h867f: y = 16'hfe00;
			16'h8680: y = 16'hfe00;
			16'h8681: y = 16'hfe00;
			16'h8682: y = 16'hfe00;
			16'h8683: y = 16'hfe00;
			16'h8684: y = 16'hfe00;
			16'h8685: y = 16'hfe00;
			16'h8686: y = 16'hfe00;
			16'h8687: y = 16'hfe00;
			16'h8688: y = 16'hfe00;
			16'h8689: y = 16'hfe00;
			16'h868a: y = 16'hfe00;
			16'h868b: y = 16'hfe00;
			16'h868c: y = 16'hfe00;
			16'h868d: y = 16'hfe00;
			16'h868e: y = 16'hfe00;
			16'h868f: y = 16'hfe00;
			16'h8690: y = 16'hfe00;
			16'h8691: y = 16'hfe00;
			16'h8692: y = 16'hfe00;
			16'h8693: y = 16'hfe00;
			16'h8694: y = 16'hfe00;
			16'h8695: y = 16'hfe00;
			16'h8696: y = 16'hfe00;
			16'h8697: y = 16'hfe00;
			16'h8698: y = 16'hfe00;
			16'h8699: y = 16'hfe00;
			16'h869a: y = 16'hfe00;
			16'h869b: y = 16'hfe00;
			16'h869c: y = 16'hfe00;
			16'h869d: y = 16'hfe00;
			16'h869e: y = 16'hfe00;
			16'h869f: y = 16'hfe00;
			16'h86a0: y = 16'hfe00;
			16'h86a1: y = 16'hfe00;
			16'h86a2: y = 16'hfe00;
			16'h86a3: y = 16'hfe00;
			16'h86a4: y = 16'hfe00;
			16'h86a5: y = 16'hfe00;
			16'h86a6: y = 16'hfe00;
			16'h86a7: y = 16'hfe00;
			16'h86a8: y = 16'hfe00;
			16'h86a9: y = 16'hfe00;
			16'h86aa: y = 16'hfe00;
			16'h86ab: y = 16'hfe00;
			16'h86ac: y = 16'hfe00;
			16'h86ad: y = 16'hfe00;
			16'h86ae: y = 16'hfe00;
			16'h86af: y = 16'hfe00;
			16'h86b0: y = 16'hfe00;
			16'h86b1: y = 16'hfe00;
			16'h86b2: y = 16'hfe00;
			16'h86b3: y = 16'hfe00;
			16'h86b4: y = 16'hfe00;
			16'h86b5: y = 16'hfe00;
			16'h86b6: y = 16'hfe00;
			16'h86b7: y = 16'hfe00;
			16'h86b8: y = 16'hfe00;
			16'h86b9: y = 16'hfe00;
			16'h86ba: y = 16'hfe00;
			16'h86bb: y = 16'hfe00;
			16'h86bc: y = 16'hfe00;
			16'h86bd: y = 16'hfe00;
			16'h86be: y = 16'hfe00;
			16'h86bf: y = 16'hfe00;
			16'h86c0: y = 16'hfe00;
			16'h86c1: y = 16'hfe00;
			16'h86c2: y = 16'hfe00;
			16'h86c3: y = 16'hfe00;
			16'h86c4: y = 16'hfe00;
			16'h86c5: y = 16'hfe00;
			16'h86c6: y = 16'hfe00;
			16'h86c7: y = 16'hfe00;
			16'h86c8: y = 16'hfe00;
			16'h86c9: y = 16'hfe00;
			16'h86ca: y = 16'hfe00;
			16'h86cb: y = 16'hfe00;
			16'h86cc: y = 16'hfe00;
			16'h86cd: y = 16'hfe00;
			16'h86ce: y = 16'hfe00;
			16'h86cf: y = 16'hfe00;
			16'h86d0: y = 16'hfe00;
			16'h86d1: y = 16'hfe00;
			16'h86d2: y = 16'hfe00;
			16'h86d3: y = 16'hfe00;
			16'h86d4: y = 16'hfe00;
			16'h86d5: y = 16'hfe00;
			16'h86d6: y = 16'hfe00;
			16'h86d7: y = 16'hfe00;
			16'h86d8: y = 16'hfe00;
			16'h86d9: y = 16'hfe00;
			16'h86da: y = 16'hfe00;
			16'h86db: y = 16'hfe00;
			16'h86dc: y = 16'hfe00;
			16'h86dd: y = 16'hfe00;
			16'h86de: y = 16'hfe00;
			16'h86df: y = 16'hfe00;
			16'h86e0: y = 16'hfe00;
			16'h86e1: y = 16'hfe00;
			16'h86e2: y = 16'hfe00;
			16'h86e3: y = 16'hfe00;
			16'h86e4: y = 16'hfe00;
			16'h86e5: y = 16'hfe00;
			16'h86e6: y = 16'hfe00;
			16'h86e7: y = 16'hfe00;
			16'h86e8: y = 16'hfe00;
			16'h86e9: y = 16'hfe00;
			16'h86ea: y = 16'hfe00;
			16'h86eb: y = 16'hfe00;
			16'h86ec: y = 16'hfe00;
			16'h86ed: y = 16'hfe00;
			16'h86ee: y = 16'hfe00;
			16'h86ef: y = 16'hfe00;
			16'h86f0: y = 16'hfe00;
			16'h86f1: y = 16'hfe00;
			16'h86f2: y = 16'hfe00;
			16'h86f3: y = 16'hfe00;
			16'h86f4: y = 16'hfe00;
			16'h86f5: y = 16'hfe00;
			16'h86f6: y = 16'hfe00;
			16'h86f7: y = 16'hfe00;
			16'h86f8: y = 16'hfe00;
			16'h86f9: y = 16'hfe00;
			16'h86fa: y = 16'hfe00;
			16'h86fb: y = 16'hfe00;
			16'h86fc: y = 16'hfe00;
			16'h86fd: y = 16'hfe00;
			16'h86fe: y = 16'hfe00;
			16'h86ff: y = 16'hfe00;
			16'h8700: y = 16'hfe00;
			16'h8701: y = 16'hfe00;
			16'h8702: y = 16'hfe00;
			16'h8703: y = 16'hfe00;
			16'h8704: y = 16'hfe00;
			16'h8705: y = 16'hfe00;
			16'h8706: y = 16'hfe00;
			16'h8707: y = 16'hfe00;
			16'h8708: y = 16'hfe00;
			16'h8709: y = 16'hfe00;
			16'h870a: y = 16'hfe00;
			16'h870b: y = 16'hfe00;
			16'h870c: y = 16'hfe00;
			16'h870d: y = 16'hfe00;
			16'h870e: y = 16'hfe00;
			16'h870f: y = 16'hfe00;
			16'h8710: y = 16'hfe00;
			16'h8711: y = 16'hfe00;
			16'h8712: y = 16'hfe00;
			16'h8713: y = 16'hfe00;
			16'h8714: y = 16'hfe00;
			16'h8715: y = 16'hfe00;
			16'h8716: y = 16'hfe00;
			16'h8717: y = 16'hfe00;
			16'h8718: y = 16'hfe00;
			16'h8719: y = 16'hfe00;
			16'h871a: y = 16'hfe00;
			16'h871b: y = 16'hfe00;
			16'h871c: y = 16'hfe00;
			16'h871d: y = 16'hfe00;
			16'h871e: y = 16'hfe00;
			16'h871f: y = 16'hfe00;
			16'h8720: y = 16'hfe00;
			16'h8721: y = 16'hfe00;
			16'h8722: y = 16'hfe00;
			16'h8723: y = 16'hfe00;
			16'h8724: y = 16'hfe00;
			16'h8725: y = 16'hfe00;
			16'h8726: y = 16'hfe00;
			16'h8727: y = 16'hfe00;
			16'h8728: y = 16'hfe00;
			16'h8729: y = 16'hfe00;
			16'h872a: y = 16'hfe00;
			16'h872b: y = 16'hfe00;
			16'h872c: y = 16'hfe00;
			16'h872d: y = 16'hfe00;
			16'h872e: y = 16'hfe00;
			16'h872f: y = 16'hfe00;
			16'h8730: y = 16'hfe00;
			16'h8731: y = 16'hfe00;
			16'h8732: y = 16'hfe00;
			16'h8733: y = 16'hfe00;
			16'h8734: y = 16'hfe00;
			16'h8735: y = 16'hfe00;
			16'h8736: y = 16'hfe00;
			16'h8737: y = 16'hfe00;
			16'h8738: y = 16'hfe00;
			16'h8739: y = 16'hfe00;
			16'h873a: y = 16'hfe00;
			16'h873b: y = 16'hfe00;
			16'h873c: y = 16'hfe00;
			16'h873d: y = 16'hfe00;
			16'h873e: y = 16'hfe00;
			16'h873f: y = 16'hfe00;
			16'h8740: y = 16'hfe00;
			16'h8741: y = 16'hfe00;
			16'h8742: y = 16'hfe00;
			16'h8743: y = 16'hfe00;
			16'h8744: y = 16'hfe00;
			16'h8745: y = 16'hfe00;
			16'h8746: y = 16'hfe00;
			16'h8747: y = 16'hfe00;
			16'h8748: y = 16'hfe00;
			16'h8749: y = 16'hfe00;
			16'h874a: y = 16'hfe00;
			16'h874b: y = 16'hfe00;
			16'h874c: y = 16'hfe00;
			16'h874d: y = 16'hfe00;
			16'h874e: y = 16'hfe00;
			16'h874f: y = 16'hfe00;
			16'h8750: y = 16'hfe00;
			16'h8751: y = 16'hfe00;
			16'h8752: y = 16'hfe00;
			16'h8753: y = 16'hfe00;
			16'h8754: y = 16'hfe00;
			16'h8755: y = 16'hfe00;
			16'h8756: y = 16'hfe00;
			16'h8757: y = 16'hfe00;
			16'h8758: y = 16'hfe00;
			16'h8759: y = 16'hfe00;
			16'h875a: y = 16'hfe00;
			16'h875b: y = 16'hfe00;
			16'h875c: y = 16'hfe00;
			16'h875d: y = 16'hfe00;
			16'h875e: y = 16'hfe00;
			16'h875f: y = 16'hfe00;
			16'h8760: y = 16'hfe00;
			16'h8761: y = 16'hfe00;
			16'h8762: y = 16'hfe00;
			16'h8763: y = 16'hfe00;
			16'h8764: y = 16'hfe00;
			16'h8765: y = 16'hfe00;
			16'h8766: y = 16'hfe00;
			16'h8767: y = 16'hfe00;
			16'h8768: y = 16'hfe00;
			16'h8769: y = 16'hfe00;
			16'h876a: y = 16'hfe00;
			16'h876b: y = 16'hfe00;
			16'h876c: y = 16'hfe00;
			16'h876d: y = 16'hfe00;
			16'h876e: y = 16'hfe00;
			16'h876f: y = 16'hfe00;
			16'h8770: y = 16'hfe00;
			16'h8771: y = 16'hfe00;
			16'h8772: y = 16'hfe00;
			16'h8773: y = 16'hfe00;
			16'h8774: y = 16'hfe00;
			16'h8775: y = 16'hfe00;
			16'h8776: y = 16'hfe00;
			16'h8777: y = 16'hfe00;
			16'h8778: y = 16'hfe00;
			16'h8779: y = 16'hfe00;
			16'h877a: y = 16'hfe00;
			16'h877b: y = 16'hfe00;
			16'h877c: y = 16'hfe00;
			16'h877d: y = 16'hfe00;
			16'h877e: y = 16'hfe00;
			16'h877f: y = 16'hfe00;
			16'h8780: y = 16'hfe00;
			16'h8781: y = 16'hfe00;
			16'h8782: y = 16'hfe00;
			16'h8783: y = 16'hfe00;
			16'h8784: y = 16'hfe00;
			16'h8785: y = 16'hfe00;
			16'h8786: y = 16'hfe00;
			16'h8787: y = 16'hfe00;
			16'h8788: y = 16'hfe00;
			16'h8789: y = 16'hfe00;
			16'h878a: y = 16'hfe00;
			16'h878b: y = 16'hfe00;
			16'h878c: y = 16'hfe00;
			16'h878d: y = 16'hfe00;
			16'h878e: y = 16'hfe00;
			16'h878f: y = 16'hfe00;
			16'h8790: y = 16'hfe00;
			16'h8791: y = 16'hfe00;
			16'h8792: y = 16'hfe00;
			16'h8793: y = 16'hfe00;
			16'h8794: y = 16'hfe00;
			16'h8795: y = 16'hfe00;
			16'h8796: y = 16'hfe00;
			16'h8797: y = 16'hfe00;
			16'h8798: y = 16'hfe00;
			16'h8799: y = 16'hfe00;
			16'h879a: y = 16'hfe00;
			16'h879b: y = 16'hfe00;
			16'h879c: y = 16'hfe00;
			16'h879d: y = 16'hfe00;
			16'h879e: y = 16'hfe00;
			16'h879f: y = 16'hfe00;
			16'h87a0: y = 16'hfe00;
			16'h87a1: y = 16'hfe00;
			16'h87a2: y = 16'hfe00;
			16'h87a3: y = 16'hfe00;
			16'h87a4: y = 16'hfe00;
			16'h87a5: y = 16'hfe00;
			16'h87a6: y = 16'hfe00;
			16'h87a7: y = 16'hfe00;
			16'h87a8: y = 16'hfe00;
			16'h87a9: y = 16'hfe00;
			16'h87aa: y = 16'hfe00;
			16'h87ab: y = 16'hfe00;
			16'h87ac: y = 16'hfe00;
			16'h87ad: y = 16'hfe00;
			16'h87ae: y = 16'hfe00;
			16'h87af: y = 16'hfe00;
			16'h87b0: y = 16'hfe00;
			16'h87b1: y = 16'hfe00;
			16'h87b2: y = 16'hfe00;
			16'h87b3: y = 16'hfe00;
			16'h87b4: y = 16'hfe00;
			16'h87b5: y = 16'hfe00;
			16'h87b6: y = 16'hfe00;
			16'h87b7: y = 16'hfe00;
			16'h87b8: y = 16'hfe00;
			16'h87b9: y = 16'hfe00;
			16'h87ba: y = 16'hfe00;
			16'h87bb: y = 16'hfe00;
			16'h87bc: y = 16'hfe00;
			16'h87bd: y = 16'hfe00;
			16'h87be: y = 16'hfe00;
			16'h87bf: y = 16'hfe00;
			16'h87c0: y = 16'hfe00;
			16'h87c1: y = 16'hfe00;
			16'h87c2: y = 16'hfe00;
			16'h87c3: y = 16'hfe00;
			16'h87c4: y = 16'hfe00;
			16'h87c5: y = 16'hfe00;
			16'h87c6: y = 16'hfe00;
			16'h87c7: y = 16'hfe00;
			16'h87c8: y = 16'hfe00;
			16'h87c9: y = 16'hfe00;
			16'h87ca: y = 16'hfe00;
			16'h87cb: y = 16'hfe00;
			16'h87cc: y = 16'hfe00;
			16'h87cd: y = 16'hfe00;
			16'h87ce: y = 16'hfe00;
			16'h87cf: y = 16'hfe00;
			16'h87d0: y = 16'hfe00;
			16'h87d1: y = 16'hfe00;
			16'h87d2: y = 16'hfe00;
			16'h87d3: y = 16'hfe00;
			16'h87d4: y = 16'hfe00;
			16'h87d5: y = 16'hfe00;
			16'h87d6: y = 16'hfe00;
			16'h87d7: y = 16'hfe00;
			16'h87d8: y = 16'hfe00;
			16'h87d9: y = 16'hfe00;
			16'h87da: y = 16'hfe00;
			16'h87db: y = 16'hfe00;
			16'h87dc: y = 16'hfe00;
			16'h87dd: y = 16'hfe00;
			16'h87de: y = 16'hfe00;
			16'h87df: y = 16'hfe00;
			16'h87e0: y = 16'hfe00;
			16'h87e1: y = 16'hfe00;
			16'h87e2: y = 16'hfe00;
			16'h87e3: y = 16'hfe00;
			16'h87e4: y = 16'hfe00;
			16'h87e5: y = 16'hfe00;
			16'h87e6: y = 16'hfe00;
			16'h87e7: y = 16'hfe00;
			16'h87e8: y = 16'hfe00;
			16'h87e9: y = 16'hfe00;
			16'h87ea: y = 16'hfe00;
			16'h87eb: y = 16'hfe00;
			16'h87ec: y = 16'hfe00;
			16'h87ed: y = 16'hfe00;
			16'h87ee: y = 16'hfe00;
			16'h87ef: y = 16'hfe00;
			16'h87f0: y = 16'hfe00;
			16'h87f1: y = 16'hfe00;
			16'h87f2: y = 16'hfe00;
			16'h87f3: y = 16'hfe00;
			16'h87f4: y = 16'hfe00;
			16'h87f5: y = 16'hfe00;
			16'h87f6: y = 16'hfe00;
			16'h87f7: y = 16'hfe00;
			16'h87f8: y = 16'hfe00;
			16'h87f9: y = 16'hfe00;
			16'h87fa: y = 16'hfe00;
			16'h87fb: y = 16'hfe00;
			16'h87fc: y = 16'hfe00;
			16'h87fd: y = 16'hfe00;
			16'h87fe: y = 16'hfe00;
			16'h87ff: y = 16'hfe00;
			16'h8800: y = 16'hfe00;
			16'h8801: y = 16'hfe00;
			16'h8802: y = 16'hfe00;
			16'h8803: y = 16'hfe00;
			16'h8804: y = 16'hfe00;
			16'h8805: y = 16'hfe00;
			16'h8806: y = 16'hfe00;
			16'h8807: y = 16'hfe00;
			16'h8808: y = 16'hfe00;
			16'h8809: y = 16'hfe00;
			16'h880a: y = 16'hfe00;
			16'h880b: y = 16'hfe00;
			16'h880c: y = 16'hfe00;
			16'h880d: y = 16'hfe00;
			16'h880e: y = 16'hfe00;
			16'h880f: y = 16'hfe00;
			16'h8810: y = 16'hfe00;
			16'h8811: y = 16'hfe00;
			16'h8812: y = 16'hfe00;
			16'h8813: y = 16'hfe00;
			16'h8814: y = 16'hfe00;
			16'h8815: y = 16'hfe00;
			16'h8816: y = 16'hfe00;
			16'h8817: y = 16'hfe00;
			16'h8818: y = 16'hfe00;
			16'h8819: y = 16'hfe00;
			16'h881a: y = 16'hfe00;
			16'h881b: y = 16'hfe00;
			16'h881c: y = 16'hfe00;
			16'h881d: y = 16'hfe00;
			16'h881e: y = 16'hfe00;
			16'h881f: y = 16'hfe00;
			16'h8820: y = 16'hfe00;
			16'h8821: y = 16'hfe00;
			16'h8822: y = 16'hfe00;
			16'h8823: y = 16'hfe00;
			16'h8824: y = 16'hfe00;
			16'h8825: y = 16'hfe00;
			16'h8826: y = 16'hfe00;
			16'h8827: y = 16'hfe00;
			16'h8828: y = 16'hfe00;
			16'h8829: y = 16'hfe00;
			16'h882a: y = 16'hfe00;
			16'h882b: y = 16'hfe00;
			16'h882c: y = 16'hfe00;
			16'h882d: y = 16'hfe00;
			16'h882e: y = 16'hfe00;
			16'h882f: y = 16'hfe00;
			16'h8830: y = 16'hfe00;
			16'h8831: y = 16'hfe00;
			16'h8832: y = 16'hfe00;
			16'h8833: y = 16'hfe00;
			16'h8834: y = 16'hfe00;
			16'h8835: y = 16'hfe00;
			16'h8836: y = 16'hfe00;
			16'h8837: y = 16'hfe00;
			16'h8838: y = 16'hfe00;
			16'h8839: y = 16'hfe00;
			16'h883a: y = 16'hfe00;
			16'h883b: y = 16'hfe00;
			16'h883c: y = 16'hfe00;
			16'h883d: y = 16'hfe00;
			16'h883e: y = 16'hfe00;
			16'h883f: y = 16'hfe00;
			16'h8840: y = 16'hfe00;
			16'h8841: y = 16'hfe00;
			16'h8842: y = 16'hfe00;
			16'h8843: y = 16'hfe00;
			16'h8844: y = 16'hfe00;
			16'h8845: y = 16'hfe00;
			16'h8846: y = 16'hfe00;
			16'h8847: y = 16'hfe00;
			16'h8848: y = 16'hfe00;
			16'h8849: y = 16'hfe00;
			16'h884a: y = 16'hfe00;
			16'h884b: y = 16'hfe00;
			16'h884c: y = 16'hfe00;
			16'h884d: y = 16'hfe00;
			16'h884e: y = 16'hfe00;
			16'h884f: y = 16'hfe00;
			16'h8850: y = 16'hfe00;
			16'h8851: y = 16'hfe00;
			16'h8852: y = 16'hfe00;
			16'h8853: y = 16'hfe00;
			16'h8854: y = 16'hfe00;
			16'h8855: y = 16'hfe00;
			16'h8856: y = 16'hfe00;
			16'h8857: y = 16'hfe00;
			16'h8858: y = 16'hfe00;
			16'h8859: y = 16'hfe00;
			16'h885a: y = 16'hfe00;
			16'h885b: y = 16'hfe00;
			16'h885c: y = 16'hfe00;
			16'h885d: y = 16'hfe00;
			16'h885e: y = 16'hfe00;
			16'h885f: y = 16'hfe00;
			16'h8860: y = 16'hfe00;
			16'h8861: y = 16'hfe00;
			16'h8862: y = 16'hfe00;
			16'h8863: y = 16'hfe00;
			16'h8864: y = 16'hfe00;
			16'h8865: y = 16'hfe00;
			16'h8866: y = 16'hfe00;
			16'h8867: y = 16'hfe00;
			16'h8868: y = 16'hfe00;
			16'h8869: y = 16'hfe00;
			16'h886a: y = 16'hfe00;
			16'h886b: y = 16'hfe00;
			16'h886c: y = 16'hfe00;
			16'h886d: y = 16'hfe00;
			16'h886e: y = 16'hfe00;
			16'h886f: y = 16'hfe00;
			16'h8870: y = 16'hfe00;
			16'h8871: y = 16'hfe00;
			16'h8872: y = 16'hfe00;
			16'h8873: y = 16'hfe00;
			16'h8874: y = 16'hfe00;
			16'h8875: y = 16'hfe00;
			16'h8876: y = 16'hfe00;
			16'h8877: y = 16'hfe00;
			16'h8878: y = 16'hfe00;
			16'h8879: y = 16'hfe00;
			16'h887a: y = 16'hfe00;
			16'h887b: y = 16'hfe00;
			16'h887c: y = 16'hfe00;
			16'h887d: y = 16'hfe00;
			16'h887e: y = 16'hfe00;
			16'h887f: y = 16'hfe00;
			16'h8880: y = 16'hfe00;
			16'h8881: y = 16'hfe00;
			16'h8882: y = 16'hfe00;
			16'h8883: y = 16'hfe00;
			16'h8884: y = 16'hfe00;
			16'h8885: y = 16'hfe00;
			16'h8886: y = 16'hfe00;
			16'h8887: y = 16'hfe00;
			16'h8888: y = 16'hfe00;
			16'h8889: y = 16'hfe00;
			16'h888a: y = 16'hfe00;
			16'h888b: y = 16'hfe00;
			16'h888c: y = 16'hfe00;
			16'h888d: y = 16'hfe00;
			16'h888e: y = 16'hfe00;
			16'h888f: y = 16'hfe00;
			16'h8890: y = 16'hfe00;
			16'h8891: y = 16'hfe00;
			16'h8892: y = 16'hfe00;
			16'h8893: y = 16'hfe00;
			16'h8894: y = 16'hfe00;
			16'h8895: y = 16'hfe00;
			16'h8896: y = 16'hfe00;
			16'h8897: y = 16'hfe00;
			16'h8898: y = 16'hfe00;
			16'h8899: y = 16'hfe00;
			16'h889a: y = 16'hfe00;
			16'h889b: y = 16'hfe00;
			16'h889c: y = 16'hfe00;
			16'h889d: y = 16'hfe00;
			16'h889e: y = 16'hfe00;
			16'h889f: y = 16'hfe00;
			16'h88a0: y = 16'hfe00;
			16'h88a1: y = 16'hfe00;
			16'h88a2: y = 16'hfe00;
			16'h88a3: y = 16'hfe00;
			16'h88a4: y = 16'hfe00;
			16'h88a5: y = 16'hfe00;
			16'h88a6: y = 16'hfe00;
			16'h88a7: y = 16'hfe00;
			16'h88a8: y = 16'hfe00;
			16'h88a9: y = 16'hfe00;
			16'h88aa: y = 16'hfe00;
			16'h88ab: y = 16'hfe00;
			16'h88ac: y = 16'hfe00;
			16'h88ad: y = 16'hfe00;
			16'h88ae: y = 16'hfe00;
			16'h88af: y = 16'hfe00;
			16'h88b0: y = 16'hfe00;
			16'h88b1: y = 16'hfe00;
			16'h88b2: y = 16'hfe00;
			16'h88b3: y = 16'hfe00;
			16'h88b4: y = 16'hfe00;
			16'h88b5: y = 16'hfe00;
			16'h88b6: y = 16'hfe00;
			16'h88b7: y = 16'hfe00;
			16'h88b8: y = 16'hfe00;
			16'h88b9: y = 16'hfe00;
			16'h88ba: y = 16'hfe00;
			16'h88bb: y = 16'hfe00;
			16'h88bc: y = 16'hfe00;
			16'h88bd: y = 16'hfe00;
			16'h88be: y = 16'hfe00;
			16'h88bf: y = 16'hfe00;
			16'h88c0: y = 16'hfe00;
			16'h88c1: y = 16'hfe00;
			16'h88c2: y = 16'hfe00;
			16'h88c3: y = 16'hfe00;
			16'h88c4: y = 16'hfe00;
			16'h88c5: y = 16'hfe00;
			16'h88c6: y = 16'hfe00;
			16'h88c7: y = 16'hfe00;
			16'h88c8: y = 16'hfe00;
			16'h88c9: y = 16'hfe00;
			16'h88ca: y = 16'hfe00;
			16'h88cb: y = 16'hfe00;
			16'h88cc: y = 16'hfe00;
			16'h88cd: y = 16'hfe00;
			16'h88ce: y = 16'hfe00;
			16'h88cf: y = 16'hfe00;
			16'h88d0: y = 16'hfe00;
			16'h88d1: y = 16'hfe00;
			16'h88d2: y = 16'hfe00;
			16'h88d3: y = 16'hfe00;
			16'h88d4: y = 16'hfe00;
			16'h88d5: y = 16'hfe00;
			16'h88d6: y = 16'hfe00;
			16'h88d7: y = 16'hfe00;
			16'h88d8: y = 16'hfe00;
			16'h88d9: y = 16'hfe00;
			16'h88da: y = 16'hfe00;
			16'h88db: y = 16'hfe00;
			16'h88dc: y = 16'hfe00;
			16'h88dd: y = 16'hfe00;
			16'h88de: y = 16'hfe00;
			16'h88df: y = 16'hfe00;
			16'h88e0: y = 16'hfe00;
			16'h88e1: y = 16'hfe00;
			16'h88e2: y = 16'hfe00;
			16'h88e3: y = 16'hfe00;
			16'h88e4: y = 16'hfe00;
			16'h88e5: y = 16'hfe00;
			16'h88e6: y = 16'hfe00;
			16'h88e7: y = 16'hfe00;
			16'h88e8: y = 16'hfe00;
			16'h88e9: y = 16'hfe00;
			16'h88ea: y = 16'hfe00;
			16'h88eb: y = 16'hfe00;
			16'h88ec: y = 16'hfe00;
			16'h88ed: y = 16'hfe00;
			16'h88ee: y = 16'hfe00;
			16'h88ef: y = 16'hfe00;
			16'h88f0: y = 16'hfe00;
			16'h88f1: y = 16'hfe00;
			16'h88f2: y = 16'hfe00;
			16'h88f3: y = 16'hfe00;
			16'h88f4: y = 16'hfe00;
			16'h88f5: y = 16'hfe00;
			16'h88f6: y = 16'hfe00;
			16'h88f7: y = 16'hfe00;
			16'h88f8: y = 16'hfe00;
			16'h88f9: y = 16'hfe00;
			16'h88fa: y = 16'hfe00;
			16'h88fb: y = 16'hfe00;
			16'h88fc: y = 16'hfe00;
			16'h88fd: y = 16'hfe00;
			16'h88fe: y = 16'hfe00;
			16'h88ff: y = 16'hfe00;
			16'h8900: y = 16'hfe00;
			16'h8901: y = 16'hfe00;
			16'h8902: y = 16'hfe00;
			16'h8903: y = 16'hfe00;
			16'h8904: y = 16'hfe00;
			16'h8905: y = 16'hfe00;
			16'h8906: y = 16'hfe00;
			16'h8907: y = 16'hfe00;
			16'h8908: y = 16'hfe00;
			16'h8909: y = 16'hfe00;
			16'h890a: y = 16'hfe00;
			16'h890b: y = 16'hfe00;
			16'h890c: y = 16'hfe00;
			16'h890d: y = 16'hfe00;
			16'h890e: y = 16'hfe00;
			16'h890f: y = 16'hfe00;
			16'h8910: y = 16'hfe00;
			16'h8911: y = 16'hfe00;
			16'h8912: y = 16'hfe00;
			16'h8913: y = 16'hfe00;
			16'h8914: y = 16'hfe00;
			16'h8915: y = 16'hfe00;
			16'h8916: y = 16'hfe00;
			16'h8917: y = 16'hfe00;
			16'h8918: y = 16'hfe00;
			16'h8919: y = 16'hfe00;
			16'h891a: y = 16'hfe00;
			16'h891b: y = 16'hfe00;
			16'h891c: y = 16'hfe00;
			16'h891d: y = 16'hfe00;
			16'h891e: y = 16'hfe00;
			16'h891f: y = 16'hfe00;
			16'h8920: y = 16'hfe00;
			16'h8921: y = 16'hfe00;
			16'h8922: y = 16'hfe00;
			16'h8923: y = 16'hfe00;
			16'h8924: y = 16'hfe00;
			16'h8925: y = 16'hfe00;
			16'h8926: y = 16'hfe00;
			16'h8927: y = 16'hfe00;
			16'h8928: y = 16'hfe00;
			16'h8929: y = 16'hfe00;
			16'h892a: y = 16'hfe00;
			16'h892b: y = 16'hfe00;
			16'h892c: y = 16'hfe00;
			16'h892d: y = 16'hfe00;
			16'h892e: y = 16'hfe00;
			16'h892f: y = 16'hfe00;
			16'h8930: y = 16'hfe00;
			16'h8931: y = 16'hfe00;
			16'h8932: y = 16'hfe00;
			16'h8933: y = 16'hfe00;
			16'h8934: y = 16'hfe00;
			16'h8935: y = 16'hfe00;
			16'h8936: y = 16'hfe00;
			16'h8937: y = 16'hfe00;
			16'h8938: y = 16'hfe00;
			16'h8939: y = 16'hfe00;
			16'h893a: y = 16'hfe00;
			16'h893b: y = 16'hfe00;
			16'h893c: y = 16'hfe00;
			16'h893d: y = 16'hfe00;
			16'h893e: y = 16'hfe00;
			16'h893f: y = 16'hfe00;
			16'h8940: y = 16'hfe00;
			16'h8941: y = 16'hfe00;
			16'h8942: y = 16'hfe00;
			16'h8943: y = 16'hfe00;
			16'h8944: y = 16'hfe00;
			16'h8945: y = 16'hfe00;
			16'h8946: y = 16'hfe00;
			16'h8947: y = 16'hfe00;
			16'h8948: y = 16'hfe00;
			16'h8949: y = 16'hfe00;
			16'h894a: y = 16'hfe00;
			16'h894b: y = 16'hfe00;
			16'h894c: y = 16'hfe00;
			16'h894d: y = 16'hfe00;
			16'h894e: y = 16'hfe00;
			16'h894f: y = 16'hfe00;
			16'h8950: y = 16'hfe00;
			16'h8951: y = 16'hfe00;
			16'h8952: y = 16'hfe00;
			16'h8953: y = 16'hfe00;
			16'h8954: y = 16'hfe00;
			16'h8955: y = 16'hfe00;
			16'h8956: y = 16'hfe00;
			16'h8957: y = 16'hfe00;
			16'h8958: y = 16'hfe00;
			16'h8959: y = 16'hfe00;
			16'h895a: y = 16'hfe00;
			16'h895b: y = 16'hfe00;
			16'h895c: y = 16'hfe00;
			16'h895d: y = 16'hfe00;
			16'h895e: y = 16'hfe00;
			16'h895f: y = 16'hfe00;
			16'h8960: y = 16'hfe00;
			16'h8961: y = 16'hfe00;
			16'h8962: y = 16'hfe00;
			16'h8963: y = 16'hfe00;
			16'h8964: y = 16'hfe00;
			16'h8965: y = 16'hfe00;
			16'h8966: y = 16'hfe00;
			16'h8967: y = 16'hfe00;
			16'h8968: y = 16'hfe00;
			16'h8969: y = 16'hfe00;
			16'h896a: y = 16'hfe00;
			16'h896b: y = 16'hfe00;
			16'h896c: y = 16'hfe00;
			16'h896d: y = 16'hfe00;
			16'h896e: y = 16'hfe00;
			16'h896f: y = 16'hfe00;
			16'h8970: y = 16'hfe00;
			16'h8971: y = 16'hfe00;
			16'h8972: y = 16'hfe00;
			16'h8973: y = 16'hfe00;
			16'h8974: y = 16'hfe00;
			16'h8975: y = 16'hfe00;
			16'h8976: y = 16'hfe00;
			16'h8977: y = 16'hfe00;
			16'h8978: y = 16'hfe00;
			16'h8979: y = 16'hfe00;
			16'h897a: y = 16'hfe00;
			16'h897b: y = 16'hfe00;
			16'h897c: y = 16'hfe00;
			16'h897d: y = 16'hfe00;
			16'h897e: y = 16'hfe00;
			16'h897f: y = 16'hfe00;
			16'h8980: y = 16'hfe00;
			16'h8981: y = 16'hfe00;
			16'h8982: y = 16'hfe00;
			16'h8983: y = 16'hfe00;
			16'h8984: y = 16'hfe00;
			16'h8985: y = 16'hfe00;
			16'h8986: y = 16'hfe00;
			16'h8987: y = 16'hfe00;
			16'h8988: y = 16'hfe00;
			16'h8989: y = 16'hfe00;
			16'h898a: y = 16'hfe00;
			16'h898b: y = 16'hfe00;
			16'h898c: y = 16'hfe00;
			16'h898d: y = 16'hfe00;
			16'h898e: y = 16'hfe00;
			16'h898f: y = 16'hfe00;
			16'h8990: y = 16'hfe00;
			16'h8991: y = 16'hfe00;
			16'h8992: y = 16'hfe00;
			16'h8993: y = 16'hfe00;
			16'h8994: y = 16'hfe00;
			16'h8995: y = 16'hfe00;
			16'h8996: y = 16'hfe00;
			16'h8997: y = 16'hfe00;
			16'h8998: y = 16'hfe00;
			16'h8999: y = 16'hfe00;
			16'h899a: y = 16'hfe00;
			16'h899b: y = 16'hfe00;
			16'h899c: y = 16'hfe00;
			16'h899d: y = 16'hfe00;
			16'h899e: y = 16'hfe00;
			16'h899f: y = 16'hfe00;
			16'h89a0: y = 16'hfe00;
			16'h89a1: y = 16'hfe00;
			16'h89a2: y = 16'hfe00;
			16'h89a3: y = 16'hfe00;
			16'h89a4: y = 16'hfe00;
			16'h89a5: y = 16'hfe00;
			16'h89a6: y = 16'hfe00;
			16'h89a7: y = 16'hfe00;
			16'h89a8: y = 16'hfe00;
			16'h89a9: y = 16'hfe00;
			16'h89aa: y = 16'hfe00;
			16'h89ab: y = 16'hfe00;
			16'h89ac: y = 16'hfe00;
			16'h89ad: y = 16'hfe00;
			16'h89ae: y = 16'hfe00;
			16'h89af: y = 16'hfe00;
			16'h89b0: y = 16'hfe00;
			16'h89b1: y = 16'hfe00;
			16'h89b2: y = 16'hfe00;
			16'h89b3: y = 16'hfe00;
			16'h89b4: y = 16'hfe00;
			16'h89b5: y = 16'hfe00;
			16'h89b6: y = 16'hfe00;
			16'h89b7: y = 16'hfe00;
			16'h89b8: y = 16'hfe00;
			16'h89b9: y = 16'hfe00;
			16'h89ba: y = 16'hfe00;
			16'h89bb: y = 16'hfe00;
			16'h89bc: y = 16'hfe00;
			16'h89bd: y = 16'hfe00;
			16'h89be: y = 16'hfe00;
			16'h89bf: y = 16'hfe00;
			16'h89c0: y = 16'hfe00;
			16'h89c1: y = 16'hfe00;
			16'h89c2: y = 16'hfe00;
			16'h89c3: y = 16'hfe00;
			16'h89c4: y = 16'hfe00;
			16'h89c5: y = 16'hfe00;
			16'h89c6: y = 16'hfe00;
			16'h89c7: y = 16'hfe00;
			16'h89c8: y = 16'hfe00;
			16'h89c9: y = 16'hfe00;
			16'h89ca: y = 16'hfe00;
			16'h89cb: y = 16'hfe00;
			16'h89cc: y = 16'hfe00;
			16'h89cd: y = 16'hfe00;
			16'h89ce: y = 16'hfe00;
			16'h89cf: y = 16'hfe00;
			16'h89d0: y = 16'hfe00;
			16'h89d1: y = 16'hfe00;
			16'h89d2: y = 16'hfe00;
			16'h89d3: y = 16'hfe00;
			16'h89d4: y = 16'hfe00;
			16'h89d5: y = 16'hfe00;
			16'h89d6: y = 16'hfe00;
			16'h89d7: y = 16'hfe00;
			16'h89d8: y = 16'hfe00;
			16'h89d9: y = 16'hfe00;
			16'h89da: y = 16'hfe00;
			16'h89db: y = 16'hfe00;
			16'h89dc: y = 16'hfe00;
			16'h89dd: y = 16'hfe00;
			16'h89de: y = 16'hfe00;
			16'h89df: y = 16'hfe00;
			16'h89e0: y = 16'hfe00;
			16'h89e1: y = 16'hfe00;
			16'h89e2: y = 16'hfe00;
			16'h89e3: y = 16'hfe00;
			16'h89e4: y = 16'hfe00;
			16'h89e5: y = 16'hfe00;
			16'h89e6: y = 16'hfe00;
			16'h89e7: y = 16'hfe00;
			16'h89e8: y = 16'hfe00;
			16'h89e9: y = 16'hfe00;
			16'h89ea: y = 16'hfe00;
			16'h89eb: y = 16'hfe00;
			16'h89ec: y = 16'hfe00;
			16'h89ed: y = 16'hfe00;
			16'h89ee: y = 16'hfe00;
			16'h89ef: y = 16'hfe00;
			16'h89f0: y = 16'hfe00;
			16'h89f1: y = 16'hfe00;
			16'h89f2: y = 16'hfe00;
			16'h89f3: y = 16'hfe00;
			16'h89f4: y = 16'hfe00;
			16'h89f5: y = 16'hfe00;
			16'h89f6: y = 16'hfe00;
			16'h89f7: y = 16'hfe00;
			16'h89f8: y = 16'hfe00;
			16'h89f9: y = 16'hfe00;
			16'h89fa: y = 16'hfe00;
			16'h89fb: y = 16'hfe00;
			16'h89fc: y = 16'hfe00;
			16'h89fd: y = 16'hfe00;
			16'h89fe: y = 16'hfe00;
			16'h89ff: y = 16'hfe00;
			16'h8a00: y = 16'hfe00;
			16'h8a01: y = 16'hfe00;
			16'h8a02: y = 16'hfe00;
			16'h8a03: y = 16'hfe00;
			16'h8a04: y = 16'hfe00;
			16'h8a05: y = 16'hfe00;
			16'h8a06: y = 16'hfe00;
			16'h8a07: y = 16'hfe00;
			16'h8a08: y = 16'hfe00;
			16'h8a09: y = 16'hfe00;
			16'h8a0a: y = 16'hfe00;
			16'h8a0b: y = 16'hfe00;
			16'h8a0c: y = 16'hfe00;
			16'h8a0d: y = 16'hfe00;
			16'h8a0e: y = 16'hfe00;
			16'h8a0f: y = 16'hfe00;
			16'h8a10: y = 16'hfe00;
			16'h8a11: y = 16'hfe00;
			16'h8a12: y = 16'hfe00;
			16'h8a13: y = 16'hfe00;
			16'h8a14: y = 16'hfe00;
			16'h8a15: y = 16'hfe00;
			16'h8a16: y = 16'hfe00;
			16'h8a17: y = 16'hfe00;
			16'h8a18: y = 16'hfe00;
			16'h8a19: y = 16'hfe00;
			16'h8a1a: y = 16'hfe00;
			16'h8a1b: y = 16'hfe00;
			16'h8a1c: y = 16'hfe00;
			16'h8a1d: y = 16'hfe00;
			16'h8a1e: y = 16'hfe00;
			16'h8a1f: y = 16'hfe00;
			16'h8a20: y = 16'hfe00;
			16'h8a21: y = 16'hfe00;
			16'h8a22: y = 16'hfe00;
			16'h8a23: y = 16'hfe00;
			16'h8a24: y = 16'hfe00;
			16'h8a25: y = 16'hfe00;
			16'h8a26: y = 16'hfe00;
			16'h8a27: y = 16'hfe00;
			16'h8a28: y = 16'hfe00;
			16'h8a29: y = 16'hfe00;
			16'h8a2a: y = 16'hfe00;
			16'h8a2b: y = 16'hfe00;
			16'h8a2c: y = 16'hfe00;
			16'h8a2d: y = 16'hfe00;
			16'h8a2e: y = 16'hfe00;
			16'h8a2f: y = 16'hfe00;
			16'h8a30: y = 16'hfe00;
			16'h8a31: y = 16'hfe00;
			16'h8a32: y = 16'hfe00;
			16'h8a33: y = 16'hfe00;
			16'h8a34: y = 16'hfe00;
			16'h8a35: y = 16'hfe00;
			16'h8a36: y = 16'hfe00;
			16'h8a37: y = 16'hfe00;
			16'h8a38: y = 16'hfe00;
			16'h8a39: y = 16'hfe00;
			16'h8a3a: y = 16'hfe00;
			16'h8a3b: y = 16'hfe00;
			16'h8a3c: y = 16'hfe00;
			16'h8a3d: y = 16'hfe00;
			16'h8a3e: y = 16'hfe00;
			16'h8a3f: y = 16'hfe00;
			16'h8a40: y = 16'hfe00;
			16'h8a41: y = 16'hfe00;
			16'h8a42: y = 16'hfe00;
			16'h8a43: y = 16'hfe00;
			16'h8a44: y = 16'hfe00;
			16'h8a45: y = 16'hfe00;
			16'h8a46: y = 16'hfe00;
			16'h8a47: y = 16'hfe00;
			16'h8a48: y = 16'hfe00;
			16'h8a49: y = 16'hfe00;
			16'h8a4a: y = 16'hfe00;
			16'h8a4b: y = 16'hfe00;
			16'h8a4c: y = 16'hfe00;
			16'h8a4d: y = 16'hfe00;
			16'h8a4e: y = 16'hfe00;
			16'h8a4f: y = 16'hfe00;
			16'h8a50: y = 16'hfe00;
			16'h8a51: y = 16'hfe00;
			16'h8a52: y = 16'hfe00;
			16'h8a53: y = 16'hfe00;
			16'h8a54: y = 16'hfe00;
			16'h8a55: y = 16'hfe00;
			16'h8a56: y = 16'hfe00;
			16'h8a57: y = 16'hfe00;
			16'h8a58: y = 16'hfe00;
			16'h8a59: y = 16'hfe00;
			16'h8a5a: y = 16'hfe00;
			16'h8a5b: y = 16'hfe00;
			16'h8a5c: y = 16'hfe00;
			16'h8a5d: y = 16'hfe00;
			16'h8a5e: y = 16'hfe00;
			16'h8a5f: y = 16'hfe00;
			16'h8a60: y = 16'hfe00;
			16'h8a61: y = 16'hfe00;
			16'h8a62: y = 16'hfe00;
			16'h8a63: y = 16'hfe00;
			16'h8a64: y = 16'hfe00;
			16'h8a65: y = 16'hfe00;
			16'h8a66: y = 16'hfe00;
			16'h8a67: y = 16'hfe00;
			16'h8a68: y = 16'hfe00;
			16'h8a69: y = 16'hfe00;
			16'h8a6a: y = 16'hfe00;
			16'h8a6b: y = 16'hfe00;
			16'h8a6c: y = 16'hfe00;
			16'h8a6d: y = 16'hfe00;
			16'h8a6e: y = 16'hfe00;
			16'h8a6f: y = 16'hfe00;
			16'h8a70: y = 16'hfe00;
			16'h8a71: y = 16'hfe00;
			16'h8a72: y = 16'hfe00;
			16'h8a73: y = 16'hfe00;
			16'h8a74: y = 16'hfe00;
			16'h8a75: y = 16'hfe00;
			16'h8a76: y = 16'hfe00;
			16'h8a77: y = 16'hfe00;
			16'h8a78: y = 16'hfe00;
			16'h8a79: y = 16'hfe00;
			16'h8a7a: y = 16'hfe00;
			16'h8a7b: y = 16'hfe00;
			16'h8a7c: y = 16'hfe00;
			16'h8a7d: y = 16'hfe00;
			16'h8a7e: y = 16'hfe00;
			16'h8a7f: y = 16'hfe00;
			16'h8a80: y = 16'hfe00;
			16'h8a81: y = 16'hfe00;
			16'h8a82: y = 16'hfe00;
			16'h8a83: y = 16'hfe00;
			16'h8a84: y = 16'hfe00;
			16'h8a85: y = 16'hfe00;
			16'h8a86: y = 16'hfe00;
			16'h8a87: y = 16'hfe00;
			16'h8a88: y = 16'hfe00;
			16'h8a89: y = 16'hfe00;
			16'h8a8a: y = 16'hfe00;
			16'h8a8b: y = 16'hfe00;
			16'h8a8c: y = 16'hfe00;
			16'h8a8d: y = 16'hfe00;
			16'h8a8e: y = 16'hfe00;
			16'h8a8f: y = 16'hfe00;
			16'h8a90: y = 16'hfe00;
			16'h8a91: y = 16'hfe00;
			16'h8a92: y = 16'hfe00;
			16'h8a93: y = 16'hfe00;
			16'h8a94: y = 16'hfe00;
			16'h8a95: y = 16'hfe00;
			16'h8a96: y = 16'hfe00;
			16'h8a97: y = 16'hfe00;
			16'h8a98: y = 16'hfe00;
			16'h8a99: y = 16'hfe00;
			16'h8a9a: y = 16'hfe00;
			16'h8a9b: y = 16'hfe00;
			16'h8a9c: y = 16'hfe00;
			16'h8a9d: y = 16'hfe00;
			16'h8a9e: y = 16'hfe00;
			16'h8a9f: y = 16'hfe00;
			16'h8aa0: y = 16'hfe00;
			16'h8aa1: y = 16'hfe00;
			16'h8aa2: y = 16'hfe00;
			16'h8aa3: y = 16'hfe00;
			16'h8aa4: y = 16'hfe00;
			16'h8aa5: y = 16'hfe00;
			16'h8aa6: y = 16'hfe00;
			16'h8aa7: y = 16'hfe00;
			16'h8aa8: y = 16'hfe00;
			16'h8aa9: y = 16'hfe00;
			16'h8aaa: y = 16'hfe00;
			16'h8aab: y = 16'hfe00;
			16'h8aac: y = 16'hfe00;
			16'h8aad: y = 16'hfe00;
			16'h8aae: y = 16'hfe00;
			16'h8aaf: y = 16'hfe00;
			16'h8ab0: y = 16'hfe00;
			16'h8ab1: y = 16'hfe00;
			16'h8ab2: y = 16'hfe00;
			16'h8ab3: y = 16'hfe00;
			16'h8ab4: y = 16'hfe00;
			16'h8ab5: y = 16'hfe00;
			16'h8ab6: y = 16'hfe00;
			16'h8ab7: y = 16'hfe00;
			16'h8ab8: y = 16'hfe00;
			16'h8ab9: y = 16'hfe00;
			16'h8aba: y = 16'hfe00;
			16'h8abb: y = 16'hfe00;
			16'h8abc: y = 16'hfe00;
			16'h8abd: y = 16'hfe00;
			16'h8abe: y = 16'hfe00;
			16'h8abf: y = 16'hfe00;
			16'h8ac0: y = 16'hfe00;
			16'h8ac1: y = 16'hfe00;
			16'h8ac2: y = 16'hfe00;
			16'h8ac3: y = 16'hfe00;
			16'h8ac4: y = 16'hfe00;
			16'h8ac5: y = 16'hfe00;
			16'h8ac6: y = 16'hfe00;
			16'h8ac7: y = 16'hfe00;
			16'h8ac8: y = 16'hfe00;
			16'h8ac9: y = 16'hfe00;
			16'h8aca: y = 16'hfe00;
			16'h8acb: y = 16'hfe00;
			16'h8acc: y = 16'hfe00;
			16'h8acd: y = 16'hfe00;
			16'h8ace: y = 16'hfe00;
			16'h8acf: y = 16'hfe00;
			16'h8ad0: y = 16'hfe00;
			16'h8ad1: y = 16'hfe00;
			16'h8ad2: y = 16'hfe00;
			16'h8ad3: y = 16'hfe00;
			16'h8ad4: y = 16'hfe00;
			16'h8ad5: y = 16'hfe00;
			16'h8ad6: y = 16'hfe00;
			16'h8ad7: y = 16'hfe00;
			16'h8ad8: y = 16'hfe00;
			16'h8ad9: y = 16'hfe00;
			16'h8ada: y = 16'hfe00;
			16'h8adb: y = 16'hfe00;
			16'h8adc: y = 16'hfe00;
			16'h8add: y = 16'hfe00;
			16'h8ade: y = 16'hfe00;
			16'h8adf: y = 16'hfe00;
			16'h8ae0: y = 16'hfe00;
			16'h8ae1: y = 16'hfe00;
			16'h8ae2: y = 16'hfe00;
			16'h8ae3: y = 16'hfe00;
			16'h8ae4: y = 16'hfe00;
			16'h8ae5: y = 16'hfe00;
			16'h8ae6: y = 16'hfe00;
			16'h8ae7: y = 16'hfe00;
			16'h8ae8: y = 16'hfe00;
			16'h8ae9: y = 16'hfe00;
			16'h8aea: y = 16'hfe00;
			16'h8aeb: y = 16'hfe00;
			16'h8aec: y = 16'hfe00;
			16'h8aed: y = 16'hfe00;
			16'h8aee: y = 16'hfe00;
			16'h8aef: y = 16'hfe00;
			16'h8af0: y = 16'hfe00;
			16'h8af1: y = 16'hfe00;
			16'h8af2: y = 16'hfe00;
			16'h8af3: y = 16'hfe00;
			16'h8af4: y = 16'hfe00;
			16'h8af5: y = 16'hfe00;
			16'h8af6: y = 16'hfe00;
			16'h8af7: y = 16'hfe00;
			16'h8af8: y = 16'hfe00;
			16'h8af9: y = 16'hfe00;
			16'h8afa: y = 16'hfe00;
			16'h8afb: y = 16'hfe00;
			16'h8afc: y = 16'hfe00;
			16'h8afd: y = 16'hfe00;
			16'h8afe: y = 16'hfe00;
			16'h8aff: y = 16'hfe00;
			16'h8b00: y = 16'hfe00;
			16'h8b01: y = 16'hfe00;
			16'h8b02: y = 16'hfe00;
			16'h8b03: y = 16'hfe00;
			16'h8b04: y = 16'hfe00;
			16'h8b05: y = 16'hfe00;
			16'h8b06: y = 16'hfe00;
			16'h8b07: y = 16'hfe00;
			16'h8b08: y = 16'hfe00;
			16'h8b09: y = 16'hfe00;
			16'h8b0a: y = 16'hfe00;
			16'h8b0b: y = 16'hfe00;
			16'h8b0c: y = 16'hfe00;
			16'h8b0d: y = 16'hfe00;
			16'h8b0e: y = 16'hfe00;
			16'h8b0f: y = 16'hfe00;
			16'h8b10: y = 16'hfe00;
			16'h8b11: y = 16'hfe00;
			16'h8b12: y = 16'hfe00;
			16'h8b13: y = 16'hfe00;
			16'h8b14: y = 16'hfe00;
			16'h8b15: y = 16'hfe00;
			16'h8b16: y = 16'hfe00;
			16'h8b17: y = 16'hfe00;
			16'h8b18: y = 16'hfe00;
			16'h8b19: y = 16'hfe00;
			16'h8b1a: y = 16'hfe00;
			16'h8b1b: y = 16'hfe00;
			16'h8b1c: y = 16'hfe00;
			16'h8b1d: y = 16'hfe00;
			16'h8b1e: y = 16'hfe00;
			16'h8b1f: y = 16'hfe00;
			16'h8b20: y = 16'hfe00;
			16'h8b21: y = 16'hfe00;
			16'h8b22: y = 16'hfe00;
			16'h8b23: y = 16'hfe00;
			16'h8b24: y = 16'hfe00;
			16'h8b25: y = 16'hfe00;
			16'h8b26: y = 16'hfe00;
			16'h8b27: y = 16'hfe00;
			16'h8b28: y = 16'hfe00;
			16'h8b29: y = 16'hfe00;
			16'h8b2a: y = 16'hfe00;
			16'h8b2b: y = 16'hfe00;
			16'h8b2c: y = 16'hfe00;
			16'h8b2d: y = 16'hfe00;
			16'h8b2e: y = 16'hfe00;
			16'h8b2f: y = 16'hfe00;
			16'h8b30: y = 16'hfe00;
			16'h8b31: y = 16'hfe00;
			16'h8b32: y = 16'hfe00;
			16'h8b33: y = 16'hfe00;
			16'h8b34: y = 16'hfe00;
			16'h8b35: y = 16'hfe00;
			16'h8b36: y = 16'hfe00;
			16'h8b37: y = 16'hfe00;
			16'h8b38: y = 16'hfe00;
			16'h8b39: y = 16'hfe00;
			16'h8b3a: y = 16'hfe00;
			16'h8b3b: y = 16'hfe00;
			16'h8b3c: y = 16'hfe00;
			16'h8b3d: y = 16'hfe00;
			16'h8b3e: y = 16'hfe00;
			16'h8b3f: y = 16'hfe00;
			16'h8b40: y = 16'hfe00;
			16'h8b41: y = 16'hfe00;
			16'h8b42: y = 16'hfe00;
			16'h8b43: y = 16'hfe00;
			16'h8b44: y = 16'hfe00;
			16'h8b45: y = 16'hfe00;
			16'h8b46: y = 16'hfe00;
			16'h8b47: y = 16'hfe00;
			16'h8b48: y = 16'hfe00;
			16'h8b49: y = 16'hfe00;
			16'h8b4a: y = 16'hfe00;
			16'h8b4b: y = 16'hfe00;
			16'h8b4c: y = 16'hfe00;
			16'h8b4d: y = 16'hfe00;
			16'h8b4e: y = 16'hfe00;
			16'h8b4f: y = 16'hfe00;
			16'h8b50: y = 16'hfe00;
			16'h8b51: y = 16'hfe00;
			16'h8b52: y = 16'hfe00;
			16'h8b53: y = 16'hfe00;
			16'h8b54: y = 16'hfe00;
			16'h8b55: y = 16'hfe00;
			16'h8b56: y = 16'hfe00;
			16'h8b57: y = 16'hfe00;
			16'h8b58: y = 16'hfe00;
			16'h8b59: y = 16'hfe00;
			16'h8b5a: y = 16'hfe00;
			16'h8b5b: y = 16'hfe00;
			16'h8b5c: y = 16'hfe00;
			16'h8b5d: y = 16'hfe00;
			16'h8b5e: y = 16'hfe00;
			16'h8b5f: y = 16'hfe00;
			16'h8b60: y = 16'hfe00;
			16'h8b61: y = 16'hfe00;
			16'h8b62: y = 16'hfe00;
			16'h8b63: y = 16'hfe00;
			16'h8b64: y = 16'hfe00;
			16'h8b65: y = 16'hfe00;
			16'h8b66: y = 16'hfe00;
			16'h8b67: y = 16'hfe00;
			16'h8b68: y = 16'hfe00;
			16'h8b69: y = 16'hfe00;
			16'h8b6a: y = 16'hfe00;
			16'h8b6b: y = 16'hfe00;
			16'h8b6c: y = 16'hfe00;
			16'h8b6d: y = 16'hfe00;
			16'h8b6e: y = 16'hfe00;
			16'h8b6f: y = 16'hfe00;
			16'h8b70: y = 16'hfe00;
			16'h8b71: y = 16'hfe00;
			16'h8b72: y = 16'hfe00;
			16'h8b73: y = 16'hfe00;
			16'h8b74: y = 16'hfe00;
			16'h8b75: y = 16'hfe00;
			16'h8b76: y = 16'hfe00;
			16'h8b77: y = 16'hfe00;
			16'h8b78: y = 16'hfe00;
			16'h8b79: y = 16'hfe00;
			16'h8b7a: y = 16'hfe00;
			16'h8b7b: y = 16'hfe00;
			16'h8b7c: y = 16'hfe00;
			16'h8b7d: y = 16'hfe00;
			16'h8b7e: y = 16'hfe00;
			16'h8b7f: y = 16'hfe00;
			16'h8b80: y = 16'hfe00;
			16'h8b81: y = 16'hfe00;
			16'h8b82: y = 16'hfe00;
			16'h8b83: y = 16'hfe00;
			16'h8b84: y = 16'hfe00;
			16'h8b85: y = 16'hfe00;
			16'h8b86: y = 16'hfe00;
			16'h8b87: y = 16'hfe00;
			16'h8b88: y = 16'hfe00;
			16'h8b89: y = 16'hfe00;
			16'h8b8a: y = 16'hfe00;
			16'h8b8b: y = 16'hfe00;
			16'h8b8c: y = 16'hfe00;
			16'h8b8d: y = 16'hfe00;
			16'h8b8e: y = 16'hfe00;
			16'h8b8f: y = 16'hfe00;
			16'h8b90: y = 16'hfe00;
			16'h8b91: y = 16'hfe00;
			16'h8b92: y = 16'hfe00;
			16'h8b93: y = 16'hfe00;
			16'h8b94: y = 16'hfe00;
			16'h8b95: y = 16'hfe00;
			16'h8b96: y = 16'hfe00;
			16'h8b97: y = 16'hfe00;
			16'h8b98: y = 16'hfe00;
			16'h8b99: y = 16'hfe00;
			16'h8b9a: y = 16'hfe00;
			16'h8b9b: y = 16'hfe00;
			16'h8b9c: y = 16'hfe00;
			16'h8b9d: y = 16'hfe00;
			16'h8b9e: y = 16'hfe00;
			16'h8b9f: y = 16'hfe00;
			16'h8ba0: y = 16'hfe00;
			16'h8ba1: y = 16'hfe00;
			16'h8ba2: y = 16'hfe00;
			16'h8ba3: y = 16'hfe00;
			16'h8ba4: y = 16'hfe00;
			16'h8ba5: y = 16'hfe00;
			16'h8ba6: y = 16'hfe00;
			16'h8ba7: y = 16'hfe00;
			16'h8ba8: y = 16'hfe00;
			16'h8ba9: y = 16'hfe00;
			16'h8baa: y = 16'hfe00;
			16'h8bab: y = 16'hfe00;
			16'h8bac: y = 16'hfe00;
			16'h8bad: y = 16'hfe00;
			16'h8bae: y = 16'hfe00;
			16'h8baf: y = 16'hfe00;
			16'h8bb0: y = 16'hfe00;
			16'h8bb1: y = 16'hfe00;
			16'h8bb2: y = 16'hfe00;
			16'h8bb3: y = 16'hfe00;
			16'h8bb4: y = 16'hfe00;
			16'h8bb5: y = 16'hfe00;
			16'h8bb6: y = 16'hfe00;
			16'h8bb7: y = 16'hfe00;
			16'h8bb8: y = 16'hfe00;
			16'h8bb9: y = 16'hfe00;
			16'h8bba: y = 16'hfe00;
			16'h8bbb: y = 16'hfe00;
			16'h8bbc: y = 16'hfe00;
			16'h8bbd: y = 16'hfe00;
			16'h8bbe: y = 16'hfe00;
			16'h8bbf: y = 16'hfe00;
			16'h8bc0: y = 16'hfe00;
			16'h8bc1: y = 16'hfe00;
			16'h8bc2: y = 16'hfe00;
			16'h8bc3: y = 16'hfe00;
			16'h8bc4: y = 16'hfe00;
			16'h8bc5: y = 16'hfe00;
			16'h8bc6: y = 16'hfe00;
			16'h8bc7: y = 16'hfe00;
			16'h8bc8: y = 16'hfe00;
			16'h8bc9: y = 16'hfe00;
			16'h8bca: y = 16'hfe00;
			16'h8bcb: y = 16'hfe00;
			16'h8bcc: y = 16'hfe00;
			16'h8bcd: y = 16'hfe00;
			16'h8bce: y = 16'hfe00;
			16'h8bcf: y = 16'hfe00;
			16'h8bd0: y = 16'hfe00;
			16'h8bd1: y = 16'hfe00;
			16'h8bd2: y = 16'hfe00;
			16'h8bd3: y = 16'hfe00;
			16'h8bd4: y = 16'hfe00;
			16'h8bd5: y = 16'hfe00;
			16'h8bd6: y = 16'hfe00;
			16'h8bd7: y = 16'hfe00;
			16'h8bd8: y = 16'hfe00;
			16'h8bd9: y = 16'hfe00;
			16'h8bda: y = 16'hfe00;
			16'h8bdb: y = 16'hfe00;
			16'h8bdc: y = 16'hfe00;
			16'h8bdd: y = 16'hfe00;
			16'h8bde: y = 16'hfe00;
			16'h8bdf: y = 16'hfe00;
			16'h8be0: y = 16'hfe00;
			16'h8be1: y = 16'hfe00;
			16'h8be2: y = 16'hfe00;
			16'h8be3: y = 16'hfe00;
			16'h8be4: y = 16'hfe00;
			16'h8be5: y = 16'hfe00;
			16'h8be6: y = 16'hfe00;
			16'h8be7: y = 16'hfe00;
			16'h8be8: y = 16'hfe00;
			16'h8be9: y = 16'hfe00;
			16'h8bea: y = 16'hfe00;
			16'h8beb: y = 16'hfe00;
			16'h8bec: y = 16'hfe00;
			16'h8bed: y = 16'hfe00;
			16'h8bee: y = 16'hfe00;
			16'h8bef: y = 16'hfe00;
			16'h8bf0: y = 16'hfe00;
			16'h8bf1: y = 16'hfe00;
			16'h8bf2: y = 16'hfe00;
			16'h8bf3: y = 16'hfe00;
			16'h8bf4: y = 16'hfe00;
			16'h8bf5: y = 16'hfe00;
			16'h8bf6: y = 16'hfe00;
			16'h8bf7: y = 16'hfe00;
			16'h8bf8: y = 16'hfe00;
			16'h8bf9: y = 16'hfe00;
			16'h8bfa: y = 16'hfe00;
			16'h8bfb: y = 16'hfe00;
			16'h8bfc: y = 16'hfe00;
			16'h8bfd: y = 16'hfe00;
			16'h8bfe: y = 16'hfe00;
			16'h8bff: y = 16'hfe00;
			16'h8c00: y = 16'hfe00;
			16'h8c01: y = 16'hfe00;
			16'h8c02: y = 16'hfe00;
			16'h8c03: y = 16'hfe00;
			16'h8c04: y = 16'hfe00;
			16'h8c05: y = 16'hfe00;
			16'h8c06: y = 16'hfe00;
			16'h8c07: y = 16'hfe00;
			16'h8c08: y = 16'hfe00;
			16'h8c09: y = 16'hfe00;
			16'h8c0a: y = 16'hfe00;
			16'h8c0b: y = 16'hfe00;
			16'h8c0c: y = 16'hfe00;
			16'h8c0d: y = 16'hfe00;
			16'h8c0e: y = 16'hfe00;
			16'h8c0f: y = 16'hfe00;
			16'h8c10: y = 16'hfe00;
			16'h8c11: y = 16'hfe00;
			16'h8c12: y = 16'hfe00;
			16'h8c13: y = 16'hfe00;
			16'h8c14: y = 16'hfe00;
			16'h8c15: y = 16'hfe00;
			16'h8c16: y = 16'hfe00;
			16'h8c17: y = 16'hfe00;
			16'h8c18: y = 16'hfe00;
			16'h8c19: y = 16'hfe00;
			16'h8c1a: y = 16'hfe00;
			16'h8c1b: y = 16'hfe00;
			16'h8c1c: y = 16'hfe00;
			16'h8c1d: y = 16'hfe00;
			16'h8c1e: y = 16'hfe00;
			16'h8c1f: y = 16'hfe00;
			16'h8c20: y = 16'hfe00;
			16'h8c21: y = 16'hfe00;
			16'h8c22: y = 16'hfe00;
			16'h8c23: y = 16'hfe00;
			16'h8c24: y = 16'hfe00;
			16'h8c25: y = 16'hfe00;
			16'h8c26: y = 16'hfe00;
			16'h8c27: y = 16'hfe00;
			16'h8c28: y = 16'hfe00;
			16'h8c29: y = 16'hfe00;
			16'h8c2a: y = 16'hfe00;
			16'h8c2b: y = 16'hfe00;
			16'h8c2c: y = 16'hfe00;
			16'h8c2d: y = 16'hfe00;
			16'h8c2e: y = 16'hfe00;
			16'h8c2f: y = 16'hfe00;
			16'h8c30: y = 16'hfe00;
			16'h8c31: y = 16'hfe00;
			16'h8c32: y = 16'hfe00;
			16'h8c33: y = 16'hfe00;
			16'h8c34: y = 16'hfe00;
			16'h8c35: y = 16'hfe00;
			16'h8c36: y = 16'hfe00;
			16'h8c37: y = 16'hfe00;
			16'h8c38: y = 16'hfe00;
			16'h8c39: y = 16'hfe00;
			16'h8c3a: y = 16'hfe00;
			16'h8c3b: y = 16'hfe00;
			16'h8c3c: y = 16'hfe00;
			16'h8c3d: y = 16'hfe00;
			16'h8c3e: y = 16'hfe00;
			16'h8c3f: y = 16'hfe00;
			16'h8c40: y = 16'hfe00;
			16'h8c41: y = 16'hfe00;
			16'h8c42: y = 16'hfe00;
			16'h8c43: y = 16'hfe00;
			16'h8c44: y = 16'hfe00;
			16'h8c45: y = 16'hfe00;
			16'h8c46: y = 16'hfe00;
			16'h8c47: y = 16'hfe00;
			16'h8c48: y = 16'hfe00;
			16'h8c49: y = 16'hfe00;
			16'h8c4a: y = 16'hfe00;
			16'h8c4b: y = 16'hfe00;
			16'h8c4c: y = 16'hfe00;
			16'h8c4d: y = 16'hfe00;
			16'h8c4e: y = 16'hfe00;
			16'h8c4f: y = 16'hfe00;
			16'h8c50: y = 16'hfe00;
			16'h8c51: y = 16'hfe00;
			16'h8c52: y = 16'hfe00;
			16'h8c53: y = 16'hfe00;
			16'h8c54: y = 16'hfe00;
			16'h8c55: y = 16'hfe00;
			16'h8c56: y = 16'hfe00;
			16'h8c57: y = 16'hfe00;
			16'h8c58: y = 16'hfe00;
			16'h8c59: y = 16'hfe00;
			16'h8c5a: y = 16'hfe00;
			16'h8c5b: y = 16'hfe00;
			16'h8c5c: y = 16'hfe00;
			16'h8c5d: y = 16'hfe00;
			16'h8c5e: y = 16'hfe00;
			16'h8c5f: y = 16'hfe00;
			16'h8c60: y = 16'hfe00;
			16'h8c61: y = 16'hfe00;
			16'h8c62: y = 16'hfe00;
			16'h8c63: y = 16'hfe00;
			16'h8c64: y = 16'hfe00;
			16'h8c65: y = 16'hfe00;
			16'h8c66: y = 16'hfe00;
			16'h8c67: y = 16'hfe00;
			16'h8c68: y = 16'hfe00;
			16'h8c69: y = 16'hfe00;
			16'h8c6a: y = 16'hfe00;
			16'h8c6b: y = 16'hfe00;
			16'h8c6c: y = 16'hfe00;
			16'h8c6d: y = 16'hfe00;
			16'h8c6e: y = 16'hfe00;
			16'h8c6f: y = 16'hfe00;
			16'h8c70: y = 16'hfe00;
			16'h8c71: y = 16'hfe00;
			16'h8c72: y = 16'hfe00;
			16'h8c73: y = 16'hfe00;
			16'h8c74: y = 16'hfe00;
			16'h8c75: y = 16'hfe00;
			16'h8c76: y = 16'hfe00;
			16'h8c77: y = 16'hfe00;
			16'h8c78: y = 16'hfe00;
			16'h8c79: y = 16'hfe00;
			16'h8c7a: y = 16'hfe00;
			16'h8c7b: y = 16'hfe00;
			16'h8c7c: y = 16'hfe00;
			16'h8c7d: y = 16'hfe00;
			16'h8c7e: y = 16'hfe00;
			16'h8c7f: y = 16'hfe00;
			16'h8c80: y = 16'hfe00;
			16'h8c81: y = 16'hfe00;
			16'h8c82: y = 16'hfe00;
			16'h8c83: y = 16'hfe00;
			16'h8c84: y = 16'hfe00;
			16'h8c85: y = 16'hfe00;
			16'h8c86: y = 16'hfe00;
			16'h8c87: y = 16'hfe00;
			16'h8c88: y = 16'hfe00;
			16'h8c89: y = 16'hfe00;
			16'h8c8a: y = 16'hfe00;
			16'h8c8b: y = 16'hfe00;
			16'h8c8c: y = 16'hfe00;
			16'h8c8d: y = 16'hfe00;
			16'h8c8e: y = 16'hfe00;
			16'h8c8f: y = 16'hfe00;
			16'h8c90: y = 16'hfe00;
			16'h8c91: y = 16'hfe00;
			16'h8c92: y = 16'hfe00;
			16'h8c93: y = 16'hfe00;
			16'h8c94: y = 16'hfe00;
			16'h8c95: y = 16'hfe00;
			16'h8c96: y = 16'hfe00;
			16'h8c97: y = 16'hfe00;
			16'h8c98: y = 16'hfe00;
			16'h8c99: y = 16'hfe00;
			16'h8c9a: y = 16'hfe00;
			16'h8c9b: y = 16'hfe00;
			16'h8c9c: y = 16'hfe00;
			16'h8c9d: y = 16'hfe00;
			16'h8c9e: y = 16'hfe00;
			16'h8c9f: y = 16'hfe00;
			16'h8ca0: y = 16'hfe00;
			16'h8ca1: y = 16'hfe00;
			16'h8ca2: y = 16'hfe00;
			16'h8ca3: y = 16'hfe00;
			16'h8ca4: y = 16'hfe00;
			16'h8ca5: y = 16'hfe00;
			16'h8ca6: y = 16'hfe00;
			16'h8ca7: y = 16'hfe00;
			16'h8ca8: y = 16'hfe00;
			16'h8ca9: y = 16'hfe00;
			16'h8caa: y = 16'hfe00;
			16'h8cab: y = 16'hfe00;
			16'h8cac: y = 16'hfe00;
			16'h8cad: y = 16'hfe00;
			16'h8cae: y = 16'hfe00;
			16'h8caf: y = 16'hfe00;
			16'h8cb0: y = 16'hfe00;
			16'h8cb1: y = 16'hfe00;
			16'h8cb2: y = 16'hfe00;
			16'h8cb3: y = 16'hfe00;
			16'h8cb4: y = 16'hfe00;
			16'h8cb5: y = 16'hfe00;
			16'h8cb6: y = 16'hfe00;
			16'h8cb7: y = 16'hfe00;
			16'h8cb8: y = 16'hfe00;
			16'h8cb9: y = 16'hfe00;
			16'h8cba: y = 16'hfe00;
			16'h8cbb: y = 16'hfe00;
			16'h8cbc: y = 16'hfe00;
			16'h8cbd: y = 16'hfe00;
			16'h8cbe: y = 16'hfe00;
			16'h8cbf: y = 16'hfe00;
			16'h8cc0: y = 16'hfe00;
			16'h8cc1: y = 16'hfe00;
			16'h8cc2: y = 16'hfe00;
			16'h8cc3: y = 16'hfe00;
			16'h8cc4: y = 16'hfe00;
			16'h8cc5: y = 16'hfe00;
			16'h8cc6: y = 16'hfe00;
			16'h8cc7: y = 16'hfe00;
			16'h8cc8: y = 16'hfe00;
			16'h8cc9: y = 16'hfe00;
			16'h8cca: y = 16'hfe00;
			16'h8ccb: y = 16'hfe00;
			16'h8ccc: y = 16'hfe00;
			16'h8ccd: y = 16'hfe00;
			16'h8cce: y = 16'hfe00;
			16'h8ccf: y = 16'hfe00;
			16'h8cd0: y = 16'hfe00;
			16'h8cd1: y = 16'hfe00;
			16'h8cd2: y = 16'hfe00;
			16'h8cd3: y = 16'hfe00;
			16'h8cd4: y = 16'hfe00;
			16'h8cd5: y = 16'hfe00;
			16'h8cd6: y = 16'hfe00;
			16'h8cd7: y = 16'hfe00;
			16'h8cd8: y = 16'hfe00;
			16'h8cd9: y = 16'hfe00;
			16'h8cda: y = 16'hfe00;
			16'h8cdb: y = 16'hfe00;
			16'h8cdc: y = 16'hfe00;
			16'h8cdd: y = 16'hfe00;
			16'h8cde: y = 16'hfe00;
			16'h8cdf: y = 16'hfe00;
			16'h8ce0: y = 16'hfe00;
			16'h8ce1: y = 16'hfe00;
			16'h8ce2: y = 16'hfe00;
			16'h8ce3: y = 16'hfe00;
			16'h8ce4: y = 16'hfe00;
			16'h8ce5: y = 16'hfe00;
			16'h8ce6: y = 16'hfe00;
			16'h8ce7: y = 16'hfe00;
			16'h8ce8: y = 16'hfe00;
			16'h8ce9: y = 16'hfe00;
			16'h8cea: y = 16'hfe00;
			16'h8ceb: y = 16'hfe00;
			16'h8cec: y = 16'hfe00;
			16'h8ced: y = 16'hfe00;
			16'h8cee: y = 16'hfe00;
			16'h8cef: y = 16'hfe00;
			16'h8cf0: y = 16'hfe00;
			16'h8cf1: y = 16'hfe00;
			16'h8cf2: y = 16'hfe00;
			16'h8cf3: y = 16'hfe00;
			16'h8cf4: y = 16'hfe00;
			16'h8cf5: y = 16'hfe00;
			16'h8cf6: y = 16'hfe00;
			16'h8cf7: y = 16'hfe00;
			16'h8cf8: y = 16'hfe00;
			16'h8cf9: y = 16'hfe00;
			16'h8cfa: y = 16'hfe00;
			16'h8cfb: y = 16'hfe00;
			16'h8cfc: y = 16'hfe00;
			16'h8cfd: y = 16'hfe00;
			16'h8cfe: y = 16'hfe00;
			16'h8cff: y = 16'hfe00;
			16'h8d00: y = 16'hfe00;
			16'h8d01: y = 16'hfe00;
			16'h8d02: y = 16'hfe00;
			16'h8d03: y = 16'hfe00;
			16'h8d04: y = 16'hfe00;
			16'h8d05: y = 16'hfe00;
			16'h8d06: y = 16'hfe00;
			16'h8d07: y = 16'hfe00;
			16'h8d08: y = 16'hfe00;
			16'h8d09: y = 16'hfe00;
			16'h8d0a: y = 16'hfe00;
			16'h8d0b: y = 16'hfe00;
			16'h8d0c: y = 16'hfe00;
			16'h8d0d: y = 16'hfe00;
			16'h8d0e: y = 16'hfe00;
			16'h8d0f: y = 16'hfe00;
			16'h8d10: y = 16'hfe00;
			16'h8d11: y = 16'hfe00;
			16'h8d12: y = 16'hfe00;
			16'h8d13: y = 16'hfe00;
			16'h8d14: y = 16'hfe00;
			16'h8d15: y = 16'hfe00;
			16'h8d16: y = 16'hfe00;
			16'h8d17: y = 16'hfe00;
			16'h8d18: y = 16'hfe00;
			16'h8d19: y = 16'hfe00;
			16'h8d1a: y = 16'hfe00;
			16'h8d1b: y = 16'hfe00;
			16'h8d1c: y = 16'hfe00;
			16'h8d1d: y = 16'hfe00;
			16'h8d1e: y = 16'hfe00;
			16'h8d1f: y = 16'hfe00;
			16'h8d20: y = 16'hfe00;
			16'h8d21: y = 16'hfe00;
			16'h8d22: y = 16'hfe00;
			16'h8d23: y = 16'hfe00;
			16'h8d24: y = 16'hfe00;
			16'h8d25: y = 16'hfe00;
			16'h8d26: y = 16'hfe00;
			16'h8d27: y = 16'hfe00;
			16'h8d28: y = 16'hfe00;
			16'h8d29: y = 16'hfe00;
			16'h8d2a: y = 16'hfe00;
			16'h8d2b: y = 16'hfe00;
			16'h8d2c: y = 16'hfe00;
			16'h8d2d: y = 16'hfe00;
			16'h8d2e: y = 16'hfe00;
			16'h8d2f: y = 16'hfe00;
			16'h8d30: y = 16'hfe00;
			16'h8d31: y = 16'hfe00;
			16'h8d32: y = 16'hfe00;
			16'h8d33: y = 16'hfe00;
			16'h8d34: y = 16'hfe00;
			16'h8d35: y = 16'hfe00;
			16'h8d36: y = 16'hfe00;
			16'h8d37: y = 16'hfe00;
			16'h8d38: y = 16'hfe00;
			16'h8d39: y = 16'hfe00;
			16'h8d3a: y = 16'hfe00;
			16'h8d3b: y = 16'hfe00;
			16'h8d3c: y = 16'hfe00;
			16'h8d3d: y = 16'hfe00;
			16'h8d3e: y = 16'hfe00;
			16'h8d3f: y = 16'hfe00;
			16'h8d40: y = 16'hfe00;
			16'h8d41: y = 16'hfe00;
			16'h8d42: y = 16'hfe00;
			16'h8d43: y = 16'hfe00;
			16'h8d44: y = 16'hfe00;
			16'h8d45: y = 16'hfe00;
			16'h8d46: y = 16'hfe00;
			16'h8d47: y = 16'hfe00;
			16'h8d48: y = 16'hfe00;
			16'h8d49: y = 16'hfe00;
			16'h8d4a: y = 16'hfe00;
			16'h8d4b: y = 16'hfe00;
			16'h8d4c: y = 16'hfe00;
			16'h8d4d: y = 16'hfe00;
			16'h8d4e: y = 16'hfe00;
			16'h8d4f: y = 16'hfe00;
			16'h8d50: y = 16'hfe00;
			16'h8d51: y = 16'hfe00;
			16'h8d52: y = 16'hfe00;
			16'h8d53: y = 16'hfe00;
			16'h8d54: y = 16'hfe00;
			16'h8d55: y = 16'hfe00;
			16'h8d56: y = 16'hfe00;
			16'h8d57: y = 16'hfe00;
			16'h8d58: y = 16'hfe00;
			16'h8d59: y = 16'hfe00;
			16'h8d5a: y = 16'hfe00;
			16'h8d5b: y = 16'hfe00;
			16'h8d5c: y = 16'hfe00;
			16'h8d5d: y = 16'hfe00;
			16'h8d5e: y = 16'hfe00;
			16'h8d5f: y = 16'hfe00;
			16'h8d60: y = 16'hfe00;
			16'h8d61: y = 16'hfe00;
			16'h8d62: y = 16'hfe00;
			16'h8d63: y = 16'hfe00;
			16'h8d64: y = 16'hfe00;
			16'h8d65: y = 16'hfe00;
			16'h8d66: y = 16'hfe00;
			16'h8d67: y = 16'hfe00;
			16'h8d68: y = 16'hfe00;
			16'h8d69: y = 16'hfe00;
			16'h8d6a: y = 16'hfe00;
			16'h8d6b: y = 16'hfe00;
			16'h8d6c: y = 16'hfe00;
			16'h8d6d: y = 16'hfe00;
			16'h8d6e: y = 16'hfe00;
			16'h8d6f: y = 16'hfe00;
			16'h8d70: y = 16'hfe00;
			16'h8d71: y = 16'hfe00;
			16'h8d72: y = 16'hfe00;
			16'h8d73: y = 16'hfe00;
			16'h8d74: y = 16'hfe00;
			16'h8d75: y = 16'hfe00;
			16'h8d76: y = 16'hfe00;
			16'h8d77: y = 16'hfe00;
			16'h8d78: y = 16'hfe00;
			16'h8d79: y = 16'hfe00;
			16'h8d7a: y = 16'hfe00;
			16'h8d7b: y = 16'hfe00;
			16'h8d7c: y = 16'hfe00;
			16'h8d7d: y = 16'hfe00;
			16'h8d7e: y = 16'hfe00;
			16'h8d7f: y = 16'hfe00;
			16'h8d80: y = 16'hfe00;
			16'h8d81: y = 16'hfe00;
			16'h8d82: y = 16'hfe00;
			16'h8d83: y = 16'hfe00;
			16'h8d84: y = 16'hfe00;
			16'h8d85: y = 16'hfe00;
			16'h8d86: y = 16'hfe00;
			16'h8d87: y = 16'hfe00;
			16'h8d88: y = 16'hfe00;
			16'h8d89: y = 16'hfe00;
			16'h8d8a: y = 16'hfe00;
			16'h8d8b: y = 16'hfe00;
			16'h8d8c: y = 16'hfe00;
			16'h8d8d: y = 16'hfe00;
			16'h8d8e: y = 16'hfe00;
			16'h8d8f: y = 16'hfe00;
			16'h8d90: y = 16'hfe00;
			16'h8d91: y = 16'hfe00;
			16'h8d92: y = 16'hfe00;
			16'h8d93: y = 16'hfe00;
			16'h8d94: y = 16'hfe00;
			16'h8d95: y = 16'hfe00;
			16'h8d96: y = 16'hfe00;
			16'h8d97: y = 16'hfe00;
			16'h8d98: y = 16'hfe00;
			16'h8d99: y = 16'hfe00;
			16'h8d9a: y = 16'hfe00;
			16'h8d9b: y = 16'hfe00;
			16'h8d9c: y = 16'hfe00;
			16'h8d9d: y = 16'hfe00;
			16'h8d9e: y = 16'hfe00;
			16'h8d9f: y = 16'hfe00;
			16'h8da0: y = 16'hfe00;
			16'h8da1: y = 16'hfe00;
			16'h8da2: y = 16'hfe00;
			16'h8da3: y = 16'hfe00;
			16'h8da4: y = 16'hfe00;
			16'h8da5: y = 16'hfe00;
			16'h8da6: y = 16'hfe00;
			16'h8da7: y = 16'hfe00;
			16'h8da8: y = 16'hfe00;
			16'h8da9: y = 16'hfe00;
			16'h8daa: y = 16'hfe00;
			16'h8dab: y = 16'hfe00;
			16'h8dac: y = 16'hfe00;
			16'h8dad: y = 16'hfe00;
			16'h8dae: y = 16'hfe00;
			16'h8daf: y = 16'hfe00;
			16'h8db0: y = 16'hfe00;
			16'h8db1: y = 16'hfe00;
			16'h8db2: y = 16'hfe00;
			16'h8db3: y = 16'hfe00;
			16'h8db4: y = 16'hfe00;
			16'h8db5: y = 16'hfe00;
			16'h8db6: y = 16'hfe00;
			16'h8db7: y = 16'hfe00;
			16'h8db8: y = 16'hfe00;
			16'h8db9: y = 16'hfe00;
			16'h8dba: y = 16'hfe00;
			16'h8dbb: y = 16'hfe00;
			16'h8dbc: y = 16'hfe00;
			16'h8dbd: y = 16'hfe00;
			16'h8dbe: y = 16'hfe00;
			16'h8dbf: y = 16'hfe00;
			16'h8dc0: y = 16'hfe00;
			16'h8dc1: y = 16'hfe00;
			16'h8dc2: y = 16'hfe00;
			16'h8dc3: y = 16'hfe00;
			16'h8dc4: y = 16'hfe00;
			16'h8dc5: y = 16'hfe00;
			16'h8dc6: y = 16'hfe00;
			16'h8dc7: y = 16'hfe00;
			16'h8dc8: y = 16'hfe00;
			16'h8dc9: y = 16'hfe00;
			16'h8dca: y = 16'hfe00;
			16'h8dcb: y = 16'hfe00;
			16'h8dcc: y = 16'hfe00;
			16'h8dcd: y = 16'hfe00;
			16'h8dce: y = 16'hfe00;
			16'h8dcf: y = 16'hfe00;
			16'h8dd0: y = 16'hfe00;
			16'h8dd1: y = 16'hfe00;
			16'h8dd2: y = 16'hfe00;
			16'h8dd3: y = 16'hfe00;
			16'h8dd4: y = 16'hfe00;
			16'h8dd5: y = 16'hfe00;
			16'h8dd6: y = 16'hfe00;
			16'h8dd7: y = 16'hfe00;
			16'h8dd8: y = 16'hfe00;
			16'h8dd9: y = 16'hfe00;
			16'h8dda: y = 16'hfe00;
			16'h8ddb: y = 16'hfe00;
			16'h8ddc: y = 16'hfe00;
			16'h8ddd: y = 16'hfe00;
			16'h8dde: y = 16'hfe00;
			16'h8ddf: y = 16'hfe00;
			16'h8de0: y = 16'hfe00;
			16'h8de1: y = 16'hfe00;
			16'h8de2: y = 16'hfe00;
			16'h8de3: y = 16'hfe00;
			16'h8de4: y = 16'hfe00;
			16'h8de5: y = 16'hfe00;
			16'h8de6: y = 16'hfe00;
			16'h8de7: y = 16'hfe00;
			16'h8de8: y = 16'hfe00;
			16'h8de9: y = 16'hfe00;
			16'h8dea: y = 16'hfe00;
			16'h8deb: y = 16'hfe00;
			16'h8dec: y = 16'hfe00;
			16'h8ded: y = 16'hfe00;
			16'h8dee: y = 16'hfe00;
			16'h8def: y = 16'hfe00;
			16'h8df0: y = 16'hfe00;
			16'h8df1: y = 16'hfe00;
			16'h8df2: y = 16'hfe00;
			16'h8df3: y = 16'hfe00;
			16'h8df4: y = 16'hfe00;
			16'h8df5: y = 16'hfe00;
			16'h8df6: y = 16'hfe00;
			16'h8df7: y = 16'hfe00;
			16'h8df8: y = 16'hfe00;
			16'h8df9: y = 16'hfe00;
			16'h8dfa: y = 16'hfe00;
			16'h8dfb: y = 16'hfe00;
			16'h8dfc: y = 16'hfe00;
			16'h8dfd: y = 16'hfe00;
			16'h8dfe: y = 16'hfe00;
			16'h8dff: y = 16'hfe00;
			16'h8e00: y = 16'hfe00;
			16'h8e01: y = 16'hfe00;
			16'h8e02: y = 16'hfe00;
			16'h8e03: y = 16'hfe00;
			16'h8e04: y = 16'hfe00;
			16'h8e05: y = 16'hfe00;
			16'h8e06: y = 16'hfe00;
			16'h8e07: y = 16'hfe00;
			16'h8e08: y = 16'hfe00;
			16'h8e09: y = 16'hfe00;
			16'h8e0a: y = 16'hfe00;
			16'h8e0b: y = 16'hfe00;
			16'h8e0c: y = 16'hfe00;
			16'h8e0d: y = 16'hfe00;
			16'h8e0e: y = 16'hfe00;
			16'h8e0f: y = 16'hfe00;
			16'h8e10: y = 16'hfe00;
			16'h8e11: y = 16'hfe00;
			16'h8e12: y = 16'hfe00;
			16'h8e13: y = 16'hfe00;
			16'h8e14: y = 16'hfe00;
			16'h8e15: y = 16'hfe00;
			16'h8e16: y = 16'hfe00;
			16'h8e17: y = 16'hfe00;
			16'h8e18: y = 16'hfe00;
			16'h8e19: y = 16'hfe00;
			16'h8e1a: y = 16'hfe00;
			16'h8e1b: y = 16'hfe00;
			16'h8e1c: y = 16'hfe00;
			16'h8e1d: y = 16'hfe00;
			16'h8e1e: y = 16'hfe00;
			16'h8e1f: y = 16'hfe00;
			16'h8e20: y = 16'hfe00;
			16'h8e21: y = 16'hfe00;
			16'h8e22: y = 16'hfe00;
			16'h8e23: y = 16'hfe00;
			16'h8e24: y = 16'hfe00;
			16'h8e25: y = 16'hfe00;
			16'h8e26: y = 16'hfe00;
			16'h8e27: y = 16'hfe00;
			16'h8e28: y = 16'hfe00;
			16'h8e29: y = 16'hfe00;
			16'h8e2a: y = 16'hfe00;
			16'h8e2b: y = 16'hfe00;
			16'h8e2c: y = 16'hfe00;
			16'h8e2d: y = 16'hfe00;
			16'h8e2e: y = 16'hfe00;
			16'h8e2f: y = 16'hfe00;
			16'h8e30: y = 16'hfe00;
			16'h8e31: y = 16'hfe00;
			16'h8e32: y = 16'hfe00;
			16'h8e33: y = 16'hfe00;
			16'h8e34: y = 16'hfe00;
			16'h8e35: y = 16'hfe00;
			16'h8e36: y = 16'hfe00;
			16'h8e37: y = 16'hfe00;
			16'h8e38: y = 16'hfe00;
			16'h8e39: y = 16'hfe00;
			16'h8e3a: y = 16'hfe00;
			16'h8e3b: y = 16'hfe00;
			16'h8e3c: y = 16'hfe00;
			16'h8e3d: y = 16'hfe00;
			16'h8e3e: y = 16'hfe00;
			16'h8e3f: y = 16'hfe00;
			16'h8e40: y = 16'hfe00;
			16'h8e41: y = 16'hfe00;
			16'h8e42: y = 16'hfe00;
			16'h8e43: y = 16'hfe00;
			16'h8e44: y = 16'hfe00;
			16'h8e45: y = 16'hfe00;
			16'h8e46: y = 16'hfe00;
			16'h8e47: y = 16'hfe00;
			16'h8e48: y = 16'hfe00;
			16'h8e49: y = 16'hfe00;
			16'h8e4a: y = 16'hfe00;
			16'h8e4b: y = 16'hfe00;
			16'h8e4c: y = 16'hfe00;
			16'h8e4d: y = 16'hfe00;
			16'h8e4e: y = 16'hfe00;
			16'h8e4f: y = 16'hfe00;
			16'h8e50: y = 16'hfe00;
			16'h8e51: y = 16'hfe00;
			16'h8e52: y = 16'hfe00;
			16'h8e53: y = 16'hfe00;
			16'h8e54: y = 16'hfe00;
			16'h8e55: y = 16'hfe00;
			16'h8e56: y = 16'hfe00;
			16'h8e57: y = 16'hfe00;
			16'h8e58: y = 16'hfe00;
			16'h8e59: y = 16'hfe00;
			16'h8e5a: y = 16'hfe00;
			16'h8e5b: y = 16'hfe00;
			16'h8e5c: y = 16'hfe00;
			16'h8e5d: y = 16'hfe00;
			16'h8e5e: y = 16'hfe00;
			16'h8e5f: y = 16'hfe00;
			16'h8e60: y = 16'hfe00;
			16'h8e61: y = 16'hfe00;
			16'h8e62: y = 16'hfe00;
			16'h8e63: y = 16'hfe00;
			16'h8e64: y = 16'hfe00;
			16'h8e65: y = 16'hfe00;
			16'h8e66: y = 16'hfe00;
			16'h8e67: y = 16'hfe00;
			16'h8e68: y = 16'hfe00;
			16'h8e69: y = 16'hfe00;
			16'h8e6a: y = 16'hfe00;
			16'h8e6b: y = 16'hfe00;
			16'h8e6c: y = 16'hfe00;
			16'h8e6d: y = 16'hfe00;
			16'h8e6e: y = 16'hfe00;
			16'h8e6f: y = 16'hfe00;
			16'h8e70: y = 16'hfe00;
			16'h8e71: y = 16'hfe00;
			16'h8e72: y = 16'hfe00;
			16'h8e73: y = 16'hfe00;
			16'h8e74: y = 16'hfe00;
			16'h8e75: y = 16'hfe00;
			16'h8e76: y = 16'hfe00;
			16'h8e77: y = 16'hfe00;
			16'h8e78: y = 16'hfe00;
			16'h8e79: y = 16'hfe00;
			16'h8e7a: y = 16'hfe00;
			16'h8e7b: y = 16'hfe00;
			16'h8e7c: y = 16'hfe00;
			16'h8e7d: y = 16'hfe00;
			16'h8e7e: y = 16'hfe00;
			16'h8e7f: y = 16'hfe00;
			16'h8e80: y = 16'hfe00;
			16'h8e81: y = 16'hfe00;
			16'h8e82: y = 16'hfe00;
			16'h8e83: y = 16'hfe00;
			16'h8e84: y = 16'hfe00;
			16'h8e85: y = 16'hfe00;
			16'h8e86: y = 16'hfe00;
			16'h8e87: y = 16'hfe00;
			16'h8e88: y = 16'hfe00;
			16'h8e89: y = 16'hfe00;
			16'h8e8a: y = 16'hfe00;
			16'h8e8b: y = 16'hfe00;
			16'h8e8c: y = 16'hfe00;
			16'h8e8d: y = 16'hfe00;
			16'h8e8e: y = 16'hfe00;
			16'h8e8f: y = 16'hfe00;
			16'h8e90: y = 16'hfe00;
			16'h8e91: y = 16'hfe00;
			16'h8e92: y = 16'hfe00;
			16'h8e93: y = 16'hfe00;
			16'h8e94: y = 16'hfe00;
			16'h8e95: y = 16'hfe00;
			16'h8e96: y = 16'hfe00;
			16'h8e97: y = 16'hfe00;
			16'h8e98: y = 16'hfe00;
			16'h8e99: y = 16'hfe00;
			16'h8e9a: y = 16'hfe00;
			16'h8e9b: y = 16'hfe00;
			16'h8e9c: y = 16'hfe00;
			16'h8e9d: y = 16'hfe00;
			16'h8e9e: y = 16'hfe00;
			16'h8e9f: y = 16'hfe00;
			16'h8ea0: y = 16'hfe00;
			16'h8ea1: y = 16'hfe00;
			16'h8ea2: y = 16'hfe00;
			16'h8ea3: y = 16'hfe00;
			16'h8ea4: y = 16'hfe00;
			16'h8ea5: y = 16'hfe00;
			16'h8ea6: y = 16'hfe00;
			16'h8ea7: y = 16'hfe00;
			16'h8ea8: y = 16'hfe00;
			16'h8ea9: y = 16'hfe00;
			16'h8eaa: y = 16'hfe00;
			16'h8eab: y = 16'hfe00;
			16'h8eac: y = 16'hfe00;
			16'h8ead: y = 16'hfe00;
			16'h8eae: y = 16'hfe00;
			16'h8eaf: y = 16'hfe00;
			16'h8eb0: y = 16'hfe00;
			16'h8eb1: y = 16'hfe00;
			16'h8eb2: y = 16'hfe00;
			16'h8eb3: y = 16'hfe00;
			16'h8eb4: y = 16'hfe00;
			16'h8eb5: y = 16'hfe00;
			16'h8eb6: y = 16'hfe00;
			16'h8eb7: y = 16'hfe00;
			16'h8eb8: y = 16'hfe00;
			16'h8eb9: y = 16'hfe00;
			16'h8eba: y = 16'hfe00;
			16'h8ebb: y = 16'hfe00;
			16'h8ebc: y = 16'hfe00;
			16'h8ebd: y = 16'hfe00;
			16'h8ebe: y = 16'hfe00;
			16'h8ebf: y = 16'hfe00;
			16'h8ec0: y = 16'hfe00;
			16'h8ec1: y = 16'hfe00;
			16'h8ec2: y = 16'hfe00;
			16'h8ec3: y = 16'hfe00;
			16'h8ec4: y = 16'hfe00;
			16'h8ec5: y = 16'hfe00;
			16'h8ec6: y = 16'hfe00;
			16'h8ec7: y = 16'hfe00;
			16'h8ec8: y = 16'hfe00;
			16'h8ec9: y = 16'hfe00;
			16'h8eca: y = 16'hfe00;
			16'h8ecb: y = 16'hfe00;
			16'h8ecc: y = 16'hfe00;
			16'h8ecd: y = 16'hfe00;
			16'h8ece: y = 16'hfe00;
			16'h8ecf: y = 16'hfe00;
			16'h8ed0: y = 16'hfe00;
			16'h8ed1: y = 16'hfe00;
			16'h8ed2: y = 16'hfe00;
			16'h8ed3: y = 16'hfe00;
			16'h8ed4: y = 16'hfe00;
			16'h8ed5: y = 16'hfe00;
			16'h8ed6: y = 16'hfe00;
			16'h8ed7: y = 16'hfe00;
			16'h8ed8: y = 16'hfe00;
			16'h8ed9: y = 16'hfe00;
			16'h8eda: y = 16'hfe00;
			16'h8edb: y = 16'hfe00;
			16'h8edc: y = 16'hfe00;
			16'h8edd: y = 16'hfe00;
			16'h8ede: y = 16'hfe00;
			16'h8edf: y = 16'hfe00;
			16'h8ee0: y = 16'hfe00;
			16'h8ee1: y = 16'hfe00;
			16'h8ee2: y = 16'hfe00;
			16'h8ee3: y = 16'hfe00;
			16'h8ee4: y = 16'hfe00;
			16'h8ee5: y = 16'hfe00;
			16'h8ee6: y = 16'hfe00;
			16'h8ee7: y = 16'hfe00;
			16'h8ee8: y = 16'hfe00;
			16'h8ee9: y = 16'hfe00;
			16'h8eea: y = 16'hfe00;
			16'h8eeb: y = 16'hfe00;
			16'h8eec: y = 16'hfe00;
			16'h8eed: y = 16'hfe00;
			16'h8eee: y = 16'hfe00;
			16'h8eef: y = 16'hfe00;
			16'h8ef0: y = 16'hfe00;
			16'h8ef1: y = 16'hfe00;
			16'h8ef2: y = 16'hfe00;
			16'h8ef3: y = 16'hfe00;
			16'h8ef4: y = 16'hfe00;
			16'h8ef5: y = 16'hfe00;
			16'h8ef6: y = 16'hfe00;
			16'h8ef7: y = 16'hfe00;
			16'h8ef8: y = 16'hfe00;
			16'h8ef9: y = 16'hfe00;
			16'h8efa: y = 16'hfe00;
			16'h8efb: y = 16'hfe00;
			16'h8efc: y = 16'hfe00;
			16'h8efd: y = 16'hfe00;
			16'h8efe: y = 16'hfe00;
			16'h8eff: y = 16'hfe00;
			16'h8f00: y = 16'hfe00;
			16'h8f01: y = 16'hfe00;
			16'h8f02: y = 16'hfe00;
			16'h8f03: y = 16'hfe00;
			16'h8f04: y = 16'hfe00;
			16'h8f05: y = 16'hfe00;
			16'h8f06: y = 16'hfe00;
			16'h8f07: y = 16'hfe00;
			16'h8f08: y = 16'hfe00;
			16'h8f09: y = 16'hfe00;
			16'h8f0a: y = 16'hfe00;
			16'h8f0b: y = 16'hfe00;
			16'h8f0c: y = 16'hfe00;
			16'h8f0d: y = 16'hfe00;
			16'h8f0e: y = 16'hfe00;
			16'h8f0f: y = 16'hfe00;
			16'h8f10: y = 16'hfe00;
			16'h8f11: y = 16'hfe00;
			16'h8f12: y = 16'hfe00;
			16'h8f13: y = 16'hfe00;
			16'h8f14: y = 16'hfe00;
			16'h8f15: y = 16'hfe00;
			16'h8f16: y = 16'hfe00;
			16'h8f17: y = 16'hfe00;
			16'h8f18: y = 16'hfe00;
			16'h8f19: y = 16'hfe00;
			16'h8f1a: y = 16'hfe00;
			16'h8f1b: y = 16'hfe00;
			16'h8f1c: y = 16'hfe00;
			16'h8f1d: y = 16'hfe00;
			16'h8f1e: y = 16'hfe00;
			16'h8f1f: y = 16'hfe00;
			16'h8f20: y = 16'hfe00;
			16'h8f21: y = 16'hfe00;
			16'h8f22: y = 16'hfe00;
			16'h8f23: y = 16'hfe00;
			16'h8f24: y = 16'hfe00;
			16'h8f25: y = 16'hfe00;
			16'h8f26: y = 16'hfe00;
			16'h8f27: y = 16'hfe00;
			16'h8f28: y = 16'hfe00;
			16'h8f29: y = 16'hfe00;
			16'h8f2a: y = 16'hfe00;
			16'h8f2b: y = 16'hfe00;
			16'h8f2c: y = 16'hfe00;
			16'h8f2d: y = 16'hfe00;
			16'h8f2e: y = 16'hfe00;
			16'h8f2f: y = 16'hfe00;
			16'h8f30: y = 16'hfe00;
			16'h8f31: y = 16'hfe00;
			16'h8f32: y = 16'hfe00;
			16'h8f33: y = 16'hfe00;
			16'h8f34: y = 16'hfe00;
			16'h8f35: y = 16'hfe00;
			16'h8f36: y = 16'hfe00;
			16'h8f37: y = 16'hfe00;
			16'h8f38: y = 16'hfe00;
			16'h8f39: y = 16'hfe00;
			16'h8f3a: y = 16'hfe00;
			16'h8f3b: y = 16'hfe00;
			16'h8f3c: y = 16'hfe00;
			16'h8f3d: y = 16'hfe00;
			16'h8f3e: y = 16'hfe00;
			16'h8f3f: y = 16'hfe00;
			16'h8f40: y = 16'hfe00;
			16'h8f41: y = 16'hfe00;
			16'h8f42: y = 16'hfe00;
			16'h8f43: y = 16'hfe00;
			16'h8f44: y = 16'hfe00;
			16'h8f45: y = 16'hfe00;
			16'h8f46: y = 16'hfe00;
			16'h8f47: y = 16'hfe00;
			16'h8f48: y = 16'hfe00;
			16'h8f49: y = 16'hfe00;
			16'h8f4a: y = 16'hfe00;
			16'h8f4b: y = 16'hfe00;
			16'h8f4c: y = 16'hfe00;
			16'h8f4d: y = 16'hfe00;
			16'h8f4e: y = 16'hfe00;
			16'h8f4f: y = 16'hfe00;
			16'h8f50: y = 16'hfe00;
			16'h8f51: y = 16'hfe00;
			16'h8f52: y = 16'hfe00;
			16'h8f53: y = 16'hfe00;
			16'h8f54: y = 16'hfe00;
			16'h8f55: y = 16'hfe00;
			16'h8f56: y = 16'hfe00;
			16'h8f57: y = 16'hfe00;
			16'h8f58: y = 16'hfe00;
			16'h8f59: y = 16'hfe00;
			16'h8f5a: y = 16'hfe00;
			16'h8f5b: y = 16'hfe00;
			16'h8f5c: y = 16'hfe00;
			16'h8f5d: y = 16'hfe00;
			16'h8f5e: y = 16'hfe00;
			16'h8f5f: y = 16'hfe00;
			16'h8f60: y = 16'hfe00;
			16'h8f61: y = 16'hfe00;
			16'h8f62: y = 16'hfe00;
			16'h8f63: y = 16'hfe00;
			16'h8f64: y = 16'hfe00;
			16'h8f65: y = 16'hfe00;
			16'h8f66: y = 16'hfe00;
			16'h8f67: y = 16'hfe00;
			16'h8f68: y = 16'hfe00;
			16'h8f69: y = 16'hfe00;
			16'h8f6a: y = 16'hfe00;
			16'h8f6b: y = 16'hfe00;
			16'h8f6c: y = 16'hfe00;
			16'h8f6d: y = 16'hfe00;
			16'h8f6e: y = 16'hfe00;
			16'h8f6f: y = 16'hfe00;
			16'h8f70: y = 16'hfe00;
			16'h8f71: y = 16'hfe00;
			16'h8f72: y = 16'hfe00;
			16'h8f73: y = 16'hfe00;
			16'h8f74: y = 16'hfe00;
			16'h8f75: y = 16'hfe00;
			16'h8f76: y = 16'hfe00;
			16'h8f77: y = 16'hfe00;
			16'h8f78: y = 16'hfe00;
			16'h8f79: y = 16'hfe00;
			16'h8f7a: y = 16'hfe00;
			16'h8f7b: y = 16'hfe00;
			16'h8f7c: y = 16'hfe00;
			16'h8f7d: y = 16'hfe00;
			16'h8f7e: y = 16'hfe00;
			16'h8f7f: y = 16'hfe00;
			16'h8f80: y = 16'hfe00;
			16'h8f81: y = 16'hfe00;
			16'h8f82: y = 16'hfe00;
			16'h8f83: y = 16'hfe00;
			16'h8f84: y = 16'hfe00;
			16'h8f85: y = 16'hfe00;
			16'h8f86: y = 16'hfe00;
			16'h8f87: y = 16'hfe00;
			16'h8f88: y = 16'hfe00;
			16'h8f89: y = 16'hfe00;
			16'h8f8a: y = 16'hfe00;
			16'h8f8b: y = 16'hfe00;
			16'h8f8c: y = 16'hfe00;
			16'h8f8d: y = 16'hfe00;
			16'h8f8e: y = 16'hfe00;
			16'h8f8f: y = 16'hfe00;
			16'h8f90: y = 16'hfe00;
			16'h8f91: y = 16'hfe00;
			16'h8f92: y = 16'hfe00;
			16'h8f93: y = 16'hfe00;
			16'h8f94: y = 16'hfe00;
			16'h8f95: y = 16'hfe00;
			16'h8f96: y = 16'hfe00;
			16'h8f97: y = 16'hfe00;
			16'h8f98: y = 16'hfe00;
			16'h8f99: y = 16'hfe00;
			16'h8f9a: y = 16'hfe00;
			16'h8f9b: y = 16'hfe00;
			16'h8f9c: y = 16'hfe00;
			16'h8f9d: y = 16'hfe00;
			16'h8f9e: y = 16'hfe00;
			16'h8f9f: y = 16'hfe00;
			16'h8fa0: y = 16'hfe00;
			16'h8fa1: y = 16'hfe00;
			16'h8fa2: y = 16'hfe00;
			16'h8fa3: y = 16'hfe00;
			16'h8fa4: y = 16'hfe00;
			16'h8fa5: y = 16'hfe00;
			16'h8fa6: y = 16'hfe00;
			16'h8fa7: y = 16'hfe00;
			16'h8fa8: y = 16'hfe00;
			16'h8fa9: y = 16'hfe00;
			16'h8faa: y = 16'hfe00;
			16'h8fab: y = 16'hfe00;
			16'h8fac: y = 16'hfe00;
			16'h8fad: y = 16'hfe00;
			16'h8fae: y = 16'hfe00;
			16'h8faf: y = 16'hfe00;
			16'h8fb0: y = 16'hfe00;
			16'h8fb1: y = 16'hfe00;
			16'h8fb2: y = 16'hfe00;
			16'h8fb3: y = 16'hfe00;
			16'h8fb4: y = 16'hfe00;
			16'h8fb5: y = 16'hfe00;
			16'h8fb6: y = 16'hfe00;
			16'h8fb7: y = 16'hfe00;
			16'h8fb8: y = 16'hfe00;
			16'h8fb9: y = 16'hfe00;
			16'h8fba: y = 16'hfe00;
			16'h8fbb: y = 16'hfe00;
			16'h8fbc: y = 16'hfe00;
			16'h8fbd: y = 16'hfe00;
			16'h8fbe: y = 16'hfe00;
			16'h8fbf: y = 16'hfe00;
			16'h8fc0: y = 16'hfe00;
			16'h8fc1: y = 16'hfe00;
			16'h8fc2: y = 16'hfe00;
			16'h8fc3: y = 16'hfe00;
			16'h8fc4: y = 16'hfe00;
			16'h8fc5: y = 16'hfe00;
			16'h8fc6: y = 16'hfe00;
			16'h8fc7: y = 16'hfe00;
			16'h8fc8: y = 16'hfe00;
			16'h8fc9: y = 16'hfe00;
			16'h8fca: y = 16'hfe00;
			16'h8fcb: y = 16'hfe00;
			16'h8fcc: y = 16'hfe00;
			16'h8fcd: y = 16'hfe00;
			16'h8fce: y = 16'hfe00;
			16'h8fcf: y = 16'hfe00;
			16'h8fd0: y = 16'hfe00;
			16'h8fd1: y = 16'hfe00;
			16'h8fd2: y = 16'hfe00;
			16'h8fd3: y = 16'hfe00;
			16'h8fd4: y = 16'hfe00;
			16'h8fd5: y = 16'hfe00;
			16'h8fd6: y = 16'hfe00;
			16'h8fd7: y = 16'hfe00;
			16'h8fd8: y = 16'hfe00;
			16'h8fd9: y = 16'hfe00;
			16'h8fda: y = 16'hfe00;
			16'h8fdb: y = 16'hfe00;
			16'h8fdc: y = 16'hfe00;
			16'h8fdd: y = 16'hfe00;
			16'h8fde: y = 16'hfe00;
			16'h8fdf: y = 16'hfe00;
			16'h8fe0: y = 16'hfe00;
			16'h8fe1: y = 16'hfe00;
			16'h8fe2: y = 16'hfe00;
			16'h8fe3: y = 16'hfe00;
			16'h8fe4: y = 16'hfe00;
			16'h8fe5: y = 16'hfe00;
			16'h8fe6: y = 16'hfe00;
			16'h8fe7: y = 16'hfe00;
			16'h8fe8: y = 16'hfe00;
			16'h8fe9: y = 16'hfe00;
			16'h8fea: y = 16'hfe00;
			16'h8feb: y = 16'hfe00;
			16'h8fec: y = 16'hfe00;
			16'h8fed: y = 16'hfe00;
			16'h8fee: y = 16'hfe00;
			16'h8fef: y = 16'hfe00;
			16'h8ff0: y = 16'hfe00;
			16'h8ff1: y = 16'hfe00;
			16'h8ff2: y = 16'hfe00;
			16'h8ff3: y = 16'hfe00;
			16'h8ff4: y = 16'hfe00;
			16'h8ff5: y = 16'hfe00;
			16'h8ff6: y = 16'hfe00;
			16'h8ff7: y = 16'hfe00;
			16'h8ff8: y = 16'hfe00;
			16'h8ff9: y = 16'hfe00;
			16'h8ffa: y = 16'hfe00;
			16'h8ffb: y = 16'hfe00;
			16'h8ffc: y = 16'hfe00;
			16'h8ffd: y = 16'hfe00;
			16'h8ffe: y = 16'hfe00;
			16'h8fff: y = 16'hfe00;
			16'h9000: y = 16'hfe00;
			16'h9001: y = 16'hfe00;
			16'h9002: y = 16'hfe00;
			16'h9003: y = 16'hfe00;
			16'h9004: y = 16'hfe00;
			16'h9005: y = 16'hfe00;
			16'h9006: y = 16'hfe00;
			16'h9007: y = 16'hfe00;
			16'h9008: y = 16'hfe00;
			16'h9009: y = 16'hfe00;
			16'h900a: y = 16'hfe00;
			16'h900b: y = 16'hfe00;
			16'h900c: y = 16'hfe00;
			16'h900d: y = 16'hfe00;
			16'h900e: y = 16'hfe00;
			16'h900f: y = 16'hfe00;
			16'h9010: y = 16'hfe00;
			16'h9011: y = 16'hfe00;
			16'h9012: y = 16'hfe00;
			16'h9013: y = 16'hfe00;
			16'h9014: y = 16'hfe00;
			16'h9015: y = 16'hfe00;
			16'h9016: y = 16'hfe00;
			16'h9017: y = 16'hfe00;
			16'h9018: y = 16'hfe00;
			16'h9019: y = 16'hfe00;
			16'h901a: y = 16'hfe00;
			16'h901b: y = 16'hfe00;
			16'h901c: y = 16'hfe00;
			16'h901d: y = 16'hfe00;
			16'h901e: y = 16'hfe00;
			16'h901f: y = 16'hfe00;
			16'h9020: y = 16'hfe00;
			16'h9021: y = 16'hfe00;
			16'h9022: y = 16'hfe00;
			16'h9023: y = 16'hfe00;
			16'h9024: y = 16'hfe00;
			16'h9025: y = 16'hfe00;
			16'h9026: y = 16'hfe00;
			16'h9027: y = 16'hfe00;
			16'h9028: y = 16'hfe00;
			16'h9029: y = 16'hfe00;
			16'h902a: y = 16'hfe00;
			16'h902b: y = 16'hfe00;
			16'h902c: y = 16'hfe00;
			16'h902d: y = 16'hfe00;
			16'h902e: y = 16'hfe00;
			16'h902f: y = 16'hfe00;
			16'h9030: y = 16'hfe00;
			16'h9031: y = 16'hfe00;
			16'h9032: y = 16'hfe00;
			16'h9033: y = 16'hfe00;
			16'h9034: y = 16'hfe00;
			16'h9035: y = 16'hfe00;
			16'h9036: y = 16'hfe00;
			16'h9037: y = 16'hfe00;
			16'h9038: y = 16'hfe00;
			16'h9039: y = 16'hfe00;
			16'h903a: y = 16'hfe00;
			16'h903b: y = 16'hfe00;
			16'h903c: y = 16'hfe00;
			16'h903d: y = 16'hfe00;
			16'h903e: y = 16'hfe00;
			16'h903f: y = 16'hfe00;
			16'h9040: y = 16'hfe00;
			16'h9041: y = 16'hfe00;
			16'h9042: y = 16'hfe00;
			16'h9043: y = 16'hfe00;
			16'h9044: y = 16'hfe00;
			16'h9045: y = 16'hfe00;
			16'h9046: y = 16'hfe00;
			16'h9047: y = 16'hfe00;
			16'h9048: y = 16'hfe00;
			16'h9049: y = 16'hfe00;
			16'h904a: y = 16'hfe00;
			16'h904b: y = 16'hfe00;
			16'h904c: y = 16'hfe00;
			16'h904d: y = 16'hfe00;
			16'h904e: y = 16'hfe00;
			16'h904f: y = 16'hfe00;
			16'h9050: y = 16'hfe00;
			16'h9051: y = 16'hfe00;
			16'h9052: y = 16'hfe00;
			16'h9053: y = 16'hfe00;
			16'h9054: y = 16'hfe00;
			16'h9055: y = 16'hfe00;
			16'h9056: y = 16'hfe00;
			16'h9057: y = 16'hfe00;
			16'h9058: y = 16'hfe00;
			16'h9059: y = 16'hfe00;
			16'h905a: y = 16'hfe00;
			16'h905b: y = 16'hfe00;
			16'h905c: y = 16'hfe00;
			16'h905d: y = 16'hfe00;
			16'h905e: y = 16'hfe00;
			16'h905f: y = 16'hfe00;
			16'h9060: y = 16'hfe00;
			16'h9061: y = 16'hfe00;
			16'h9062: y = 16'hfe00;
			16'h9063: y = 16'hfe00;
			16'h9064: y = 16'hfe00;
			16'h9065: y = 16'hfe00;
			16'h9066: y = 16'hfe00;
			16'h9067: y = 16'hfe00;
			16'h9068: y = 16'hfe00;
			16'h9069: y = 16'hfe00;
			16'h906a: y = 16'hfe00;
			16'h906b: y = 16'hfe00;
			16'h906c: y = 16'hfe00;
			16'h906d: y = 16'hfe00;
			16'h906e: y = 16'hfe00;
			16'h906f: y = 16'hfe00;
			16'h9070: y = 16'hfe00;
			16'h9071: y = 16'hfe00;
			16'h9072: y = 16'hfe00;
			16'h9073: y = 16'hfe00;
			16'h9074: y = 16'hfe00;
			16'h9075: y = 16'hfe00;
			16'h9076: y = 16'hfe00;
			16'h9077: y = 16'hfe00;
			16'h9078: y = 16'hfe00;
			16'h9079: y = 16'hfe00;
			16'h907a: y = 16'hfe00;
			16'h907b: y = 16'hfe00;
			16'h907c: y = 16'hfe00;
			16'h907d: y = 16'hfe00;
			16'h907e: y = 16'hfe00;
			16'h907f: y = 16'hfe00;
			16'h9080: y = 16'hfe00;
			16'h9081: y = 16'hfe00;
			16'h9082: y = 16'hfe00;
			16'h9083: y = 16'hfe00;
			16'h9084: y = 16'hfe00;
			16'h9085: y = 16'hfe00;
			16'h9086: y = 16'hfe00;
			16'h9087: y = 16'hfe00;
			16'h9088: y = 16'hfe00;
			16'h9089: y = 16'hfe00;
			16'h908a: y = 16'hfe00;
			16'h908b: y = 16'hfe00;
			16'h908c: y = 16'hfe00;
			16'h908d: y = 16'hfe00;
			16'h908e: y = 16'hfe00;
			16'h908f: y = 16'hfe00;
			16'h9090: y = 16'hfe00;
			16'h9091: y = 16'hfe00;
			16'h9092: y = 16'hfe00;
			16'h9093: y = 16'hfe00;
			16'h9094: y = 16'hfe00;
			16'h9095: y = 16'hfe00;
			16'h9096: y = 16'hfe00;
			16'h9097: y = 16'hfe00;
			16'h9098: y = 16'hfe00;
			16'h9099: y = 16'hfe00;
			16'h909a: y = 16'hfe00;
			16'h909b: y = 16'hfe00;
			16'h909c: y = 16'hfe00;
			16'h909d: y = 16'hfe00;
			16'h909e: y = 16'hfe00;
			16'h909f: y = 16'hfe00;
			16'h90a0: y = 16'hfe00;
			16'h90a1: y = 16'hfe00;
			16'h90a2: y = 16'hfe00;
			16'h90a3: y = 16'hfe00;
			16'h90a4: y = 16'hfe00;
			16'h90a5: y = 16'hfe00;
			16'h90a6: y = 16'hfe00;
			16'h90a7: y = 16'hfe00;
			16'h90a8: y = 16'hfe00;
			16'h90a9: y = 16'hfe00;
			16'h90aa: y = 16'hfe00;
			16'h90ab: y = 16'hfe00;
			16'h90ac: y = 16'hfe00;
			16'h90ad: y = 16'hfe00;
			16'h90ae: y = 16'hfe00;
			16'h90af: y = 16'hfe00;
			16'h90b0: y = 16'hfe00;
			16'h90b1: y = 16'hfe00;
			16'h90b2: y = 16'hfe00;
			16'h90b3: y = 16'hfe00;
			16'h90b4: y = 16'hfe00;
			16'h90b5: y = 16'hfe00;
			16'h90b6: y = 16'hfe00;
			16'h90b7: y = 16'hfe00;
			16'h90b8: y = 16'hfe00;
			16'h90b9: y = 16'hfe00;
			16'h90ba: y = 16'hfe00;
			16'h90bb: y = 16'hfe00;
			16'h90bc: y = 16'hfe00;
			16'h90bd: y = 16'hfe00;
			16'h90be: y = 16'hfe00;
			16'h90bf: y = 16'hfe00;
			16'h90c0: y = 16'hfe00;
			16'h90c1: y = 16'hfe00;
			16'h90c2: y = 16'hfe00;
			16'h90c3: y = 16'hfe00;
			16'h90c4: y = 16'hfe00;
			16'h90c5: y = 16'hfe00;
			16'h90c6: y = 16'hfe00;
			16'h90c7: y = 16'hfe00;
			16'h90c8: y = 16'hfe00;
			16'h90c9: y = 16'hfe00;
			16'h90ca: y = 16'hfe00;
			16'h90cb: y = 16'hfe00;
			16'h90cc: y = 16'hfe00;
			16'h90cd: y = 16'hfe00;
			16'h90ce: y = 16'hfe00;
			16'h90cf: y = 16'hfe00;
			16'h90d0: y = 16'hfe00;
			16'h90d1: y = 16'hfe00;
			16'h90d2: y = 16'hfe00;
			16'h90d3: y = 16'hfe00;
			16'h90d4: y = 16'hfe00;
			16'h90d5: y = 16'hfe00;
			16'h90d6: y = 16'hfe00;
			16'h90d7: y = 16'hfe00;
			16'h90d8: y = 16'hfe00;
			16'h90d9: y = 16'hfe00;
			16'h90da: y = 16'hfe00;
			16'h90db: y = 16'hfe00;
			16'h90dc: y = 16'hfe00;
			16'h90dd: y = 16'hfe00;
			16'h90de: y = 16'hfe00;
			16'h90df: y = 16'hfe00;
			16'h90e0: y = 16'hfe00;
			16'h90e1: y = 16'hfe00;
			16'h90e2: y = 16'hfe00;
			16'h90e3: y = 16'hfe00;
			16'h90e4: y = 16'hfe00;
			16'h90e5: y = 16'hfe00;
			16'h90e6: y = 16'hfe00;
			16'h90e7: y = 16'hfe00;
			16'h90e8: y = 16'hfe00;
			16'h90e9: y = 16'hfe00;
			16'h90ea: y = 16'hfe00;
			16'h90eb: y = 16'hfe00;
			16'h90ec: y = 16'hfe00;
			16'h90ed: y = 16'hfe00;
			16'h90ee: y = 16'hfe00;
			16'h90ef: y = 16'hfe00;
			16'h90f0: y = 16'hfe00;
			16'h90f1: y = 16'hfe00;
			16'h90f2: y = 16'hfe00;
			16'h90f3: y = 16'hfe00;
			16'h90f4: y = 16'hfe00;
			16'h90f5: y = 16'hfe00;
			16'h90f6: y = 16'hfe00;
			16'h90f7: y = 16'hfe00;
			16'h90f8: y = 16'hfe00;
			16'h90f9: y = 16'hfe00;
			16'h90fa: y = 16'hfe00;
			16'h90fb: y = 16'hfe00;
			16'h90fc: y = 16'hfe00;
			16'h90fd: y = 16'hfe00;
			16'h90fe: y = 16'hfe00;
			16'h90ff: y = 16'hfe00;
			16'h9100: y = 16'hfe00;
			16'h9101: y = 16'hfe00;
			16'h9102: y = 16'hfe00;
			16'h9103: y = 16'hfe00;
			16'h9104: y = 16'hfe00;
			16'h9105: y = 16'hfe00;
			16'h9106: y = 16'hfe00;
			16'h9107: y = 16'hfe00;
			16'h9108: y = 16'hfe00;
			16'h9109: y = 16'hfe00;
			16'h910a: y = 16'hfe00;
			16'h910b: y = 16'hfe00;
			16'h910c: y = 16'hfe00;
			16'h910d: y = 16'hfe00;
			16'h910e: y = 16'hfe00;
			16'h910f: y = 16'hfe00;
			16'h9110: y = 16'hfe00;
			16'h9111: y = 16'hfe00;
			16'h9112: y = 16'hfe00;
			16'h9113: y = 16'hfe00;
			16'h9114: y = 16'hfe00;
			16'h9115: y = 16'hfe00;
			16'h9116: y = 16'hfe00;
			16'h9117: y = 16'hfe00;
			16'h9118: y = 16'hfe00;
			16'h9119: y = 16'hfe00;
			16'h911a: y = 16'hfe00;
			16'h911b: y = 16'hfe00;
			16'h911c: y = 16'hfe00;
			16'h911d: y = 16'hfe00;
			16'h911e: y = 16'hfe00;
			16'h911f: y = 16'hfe00;
			16'h9120: y = 16'hfe00;
			16'h9121: y = 16'hfe00;
			16'h9122: y = 16'hfe00;
			16'h9123: y = 16'hfe00;
			16'h9124: y = 16'hfe00;
			16'h9125: y = 16'hfe00;
			16'h9126: y = 16'hfe00;
			16'h9127: y = 16'hfe00;
			16'h9128: y = 16'hfe00;
			16'h9129: y = 16'hfe00;
			16'h912a: y = 16'hfe00;
			16'h912b: y = 16'hfe00;
			16'h912c: y = 16'hfe00;
			16'h912d: y = 16'hfe00;
			16'h912e: y = 16'hfe00;
			16'h912f: y = 16'hfe00;
			16'h9130: y = 16'hfe00;
			16'h9131: y = 16'hfe00;
			16'h9132: y = 16'hfe00;
			16'h9133: y = 16'hfe00;
			16'h9134: y = 16'hfe00;
			16'h9135: y = 16'hfe00;
			16'h9136: y = 16'hfe00;
			16'h9137: y = 16'hfe00;
			16'h9138: y = 16'hfe00;
			16'h9139: y = 16'hfe00;
			16'h913a: y = 16'hfe00;
			16'h913b: y = 16'hfe00;
			16'h913c: y = 16'hfe00;
			16'h913d: y = 16'hfe00;
			16'h913e: y = 16'hfe00;
			16'h913f: y = 16'hfe00;
			16'h9140: y = 16'hfe00;
			16'h9141: y = 16'hfe00;
			16'h9142: y = 16'hfe00;
			16'h9143: y = 16'hfe00;
			16'h9144: y = 16'hfe00;
			16'h9145: y = 16'hfe00;
			16'h9146: y = 16'hfe00;
			16'h9147: y = 16'hfe00;
			16'h9148: y = 16'hfe00;
			16'h9149: y = 16'hfe00;
			16'h914a: y = 16'hfe00;
			16'h914b: y = 16'hfe00;
			16'h914c: y = 16'hfe00;
			16'h914d: y = 16'hfe00;
			16'h914e: y = 16'hfe00;
			16'h914f: y = 16'hfe00;
			16'h9150: y = 16'hfe00;
			16'h9151: y = 16'hfe00;
			16'h9152: y = 16'hfe00;
			16'h9153: y = 16'hfe00;
			16'h9154: y = 16'hfe00;
			16'h9155: y = 16'hfe00;
			16'h9156: y = 16'hfe00;
			16'h9157: y = 16'hfe00;
			16'h9158: y = 16'hfe00;
			16'h9159: y = 16'hfe00;
			16'h915a: y = 16'hfe00;
			16'h915b: y = 16'hfe00;
			16'h915c: y = 16'hfe00;
			16'h915d: y = 16'hfe00;
			16'h915e: y = 16'hfe00;
			16'h915f: y = 16'hfe00;
			16'h9160: y = 16'hfe00;
			16'h9161: y = 16'hfe00;
			16'h9162: y = 16'hfe00;
			16'h9163: y = 16'hfe00;
			16'h9164: y = 16'hfe00;
			16'h9165: y = 16'hfe00;
			16'h9166: y = 16'hfe00;
			16'h9167: y = 16'hfe00;
			16'h9168: y = 16'hfe00;
			16'h9169: y = 16'hfe00;
			16'h916a: y = 16'hfe00;
			16'h916b: y = 16'hfe00;
			16'h916c: y = 16'hfe00;
			16'h916d: y = 16'hfe00;
			16'h916e: y = 16'hfe00;
			16'h916f: y = 16'hfe00;
			16'h9170: y = 16'hfe00;
			16'h9171: y = 16'hfe00;
			16'h9172: y = 16'hfe00;
			16'h9173: y = 16'hfe00;
			16'h9174: y = 16'hfe00;
			16'h9175: y = 16'hfe00;
			16'h9176: y = 16'hfe00;
			16'h9177: y = 16'hfe00;
			16'h9178: y = 16'hfe00;
			16'h9179: y = 16'hfe00;
			16'h917a: y = 16'hfe00;
			16'h917b: y = 16'hfe00;
			16'h917c: y = 16'hfe00;
			16'h917d: y = 16'hfe00;
			16'h917e: y = 16'hfe00;
			16'h917f: y = 16'hfe00;
			16'h9180: y = 16'hfe00;
			16'h9181: y = 16'hfe00;
			16'h9182: y = 16'hfe00;
			16'h9183: y = 16'hfe00;
			16'h9184: y = 16'hfe00;
			16'h9185: y = 16'hfe00;
			16'h9186: y = 16'hfe00;
			16'h9187: y = 16'hfe00;
			16'h9188: y = 16'hfe00;
			16'h9189: y = 16'hfe00;
			16'h918a: y = 16'hfe00;
			16'h918b: y = 16'hfe00;
			16'h918c: y = 16'hfe00;
			16'h918d: y = 16'hfe00;
			16'h918e: y = 16'hfe00;
			16'h918f: y = 16'hfe00;
			16'h9190: y = 16'hfe00;
			16'h9191: y = 16'hfe00;
			16'h9192: y = 16'hfe00;
			16'h9193: y = 16'hfe00;
			16'h9194: y = 16'hfe00;
			16'h9195: y = 16'hfe00;
			16'h9196: y = 16'hfe00;
			16'h9197: y = 16'hfe00;
			16'h9198: y = 16'hfe00;
			16'h9199: y = 16'hfe00;
			16'h919a: y = 16'hfe00;
			16'h919b: y = 16'hfe00;
			16'h919c: y = 16'hfe00;
			16'h919d: y = 16'hfe00;
			16'h919e: y = 16'hfe00;
			16'h919f: y = 16'hfe00;
			16'h91a0: y = 16'hfe00;
			16'h91a1: y = 16'hfe00;
			16'h91a2: y = 16'hfe00;
			16'h91a3: y = 16'hfe00;
			16'h91a4: y = 16'hfe00;
			16'h91a5: y = 16'hfe00;
			16'h91a6: y = 16'hfe00;
			16'h91a7: y = 16'hfe00;
			16'h91a8: y = 16'hfe00;
			16'h91a9: y = 16'hfe00;
			16'h91aa: y = 16'hfe00;
			16'h91ab: y = 16'hfe00;
			16'h91ac: y = 16'hfe00;
			16'h91ad: y = 16'hfe00;
			16'h91ae: y = 16'hfe00;
			16'h91af: y = 16'hfe00;
			16'h91b0: y = 16'hfe00;
			16'h91b1: y = 16'hfe00;
			16'h91b2: y = 16'hfe00;
			16'h91b3: y = 16'hfe00;
			16'h91b4: y = 16'hfe00;
			16'h91b5: y = 16'hfe00;
			16'h91b6: y = 16'hfe00;
			16'h91b7: y = 16'hfe00;
			16'h91b8: y = 16'hfe00;
			16'h91b9: y = 16'hfe00;
			16'h91ba: y = 16'hfe00;
			16'h91bb: y = 16'hfe00;
			16'h91bc: y = 16'hfe00;
			16'h91bd: y = 16'hfe00;
			16'h91be: y = 16'hfe00;
			16'h91bf: y = 16'hfe00;
			16'h91c0: y = 16'hfe00;
			16'h91c1: y = 16'hfe00;
			16'h91c2: y = 16'hfe00;
			16'h91c3: y = 16'hfe00;
			16'h91c4: y = 16'hfe00;
			16'h91c5: y = 16'hfe00;
			16'h91c6: y = 16'hfe00;
			16'h91c7: y = 16'hfe00;
			16'h91c8: y = 16'hfe00;
			16'h91c9: y = 16'hfe00;
			16'h91ca: y = 16'hfe00;
			16'h91cb: y = 16'hfe00;
			16'h91cc: y = 16'hfe00;
			16'h91cd: y = 16'hfe00;
			16'h91ce: y = 16'hfe00;
			16'h91cf: y = 16'hfe00;
			16'h91d0: y = 16'hfe00;
			16'h91d1: y = 16'hfe00;
			16'h91d2: y = 16'hfe00;
			16'h91d3: y = 16'hfe00;
			16'h91d4: y = 16'hfe00;
			16'h91d5: y = 16'hfe00;
			16'h91d6: y = 16'hfe00;
			16'h91d7: y = 16'hfe00;
			16'h91d8: y = 16'hfe00;
			16'h91d9: y = 16'hfe00;
			16'h91da: y = 16'hfe00;
			16'h91db: y = 16'hfe00;
			16'h91dc: y = 16'hfe00;
			16'h91dd: y = 16'hfe00;
			16'h91de: y = 16'hfe00;
			16'h91df: y = 16'hfe00;
			16'h91e0: y = 16'hfe00;
			16'h91e1: y = 16'hfe00;
			16'h91e2: y = 16'hfe00;
			16'h91e3: y = 16'hfe00;
			16'h91e4: y = 16'hfe00;
			16'h91e5: y = 16'hfe00;
			16'h91e6: y = 16'hfe00;
			16'h91e7: y = 16'hfe00;
			16'h91e8: y = 16'hfe00;
			16'h91e9: y = 16'hfe00;
			16'h91ea: y = 16'hfe00;
			16'h91eb: y = 16'hfe00;
			16'h91ec: y = 16'hfe00;
			16'h91ed: y = 16'hfe00;
			16'h91ee: y = 16'hfe00;
			16'h91ef: y = 16'hfe00;
			16'h91f0: y = 16'hfe00;
			16'h91f1: y = 16'hfe00;
			16'h91f2: y = 16'hfe00;
			16'h91f3: y = 16'hfe00;
			16'h91f4: y = 16'hfe00;
			16'h91f5: y = 16'hfe00;
			16'h91f6: y = 16'hfe00;
			16'h91f7: y = 16'hfe00;
			16'h91f8: y = 16'hfe00;
			16'h91f9: y = 16'hfe00;
			16'h91fa: y = 16'hfe00;
			16'h91fb: y = 16'hfe00;
			16'h91fc: y = 16'hfe00;
			16'h91fd: y = 16'hfe00;
			16'h91fe: y = 16'hfe00;
			16'h91ff: y = 16'hfe00;
			16'h9200: y = 16'hfe00;
			16'h9201: y = 16'hfe00;
			16'h9202: y = 16'hfe00;
			16'h9203: y = 16'hfe00;
			16'h9204: y = 16'hfe00;
			16'h9205: y = 16'hfe00;
			16'h9206: y = 16'hfe00;
			16'h9207: y = 16'hfe00;
			16'h9208: y = 16'hfe00;
			16'h9209: y = 16'hfe00;
			16'h920a: y = 16'hfe00;
			16'h920b: y = 16'hfe00;
			16'h920c: y = 16'hfe00;
			16'h920d: y = 16'hfe00;
			16'h920e: y = 16'hfe00;
			16'h920f: y = 16'hfe00;
			16'h9210: y = 16'hfe00;
			16'h9211: y = 16'hfe00;
			16'h9212: y = 16'hfe00;
			16'h9213: y = 16'hfe00;
			16'h9214: y = 16'hfe00;
			16'h9215: y = 16'hfe00;
			16'h9216: y = 16'hfe00;
			16'h9217: y = 16'hfe00;
			16'h9218: y = 16'hfe00;
			16'h9219: y = 16'hfe00;
			16'h921a: y = 16'hfe00;
			16'h921b: y = 16'hfe00;
			16'h921c: y = 16'hfe00;
			16'h921d: y = 16'hfe00;
			16'h921e: y = 16'hfe00;
			16'h921f: y = 16'hfe00;
			16'h9220: y = 16'hfe00;
			16'h9221: y = 16'hfe00;
			16'h9222: y = 16'hfe00;
			16'h9223: y = 16'hfe00;
			16'h9224: y = 16'hfe00;
			16'h9225: y = 16'hfe00;
			16'h9226: y = 16'hfe00;
			16'h9227: y = 16'hfe00;
			16'h9228: y = 16'hfe00;
			16'h9229: y = 16'hfe00;
			16'h922a: y = 16'hfe00;
			16'h922b: y = 16'hfe00;
			16'h922c: y = 16'hfe00;
			16'h922d: y = 16'hfe00;
			16'h922e: y = 16'hfe00;
			16'h922f: y = 16'hfe00;
			16'h9230: y = 16'hfe00;
			16'h9231: y = 16'hfe00;
			16'h9232: y = 16'hfe00;
			16'h9233: y = 16'hfe00;
			16'h9234: y = 16'hfe00;
			16'h9235: y = 16'hfe00;
			16'h9236: y = 16'hfe00;
			16'h9237: y = 16'hfe00;
			16'h9238: y = 16'hfe00;
			16'h9239: y = 16'hfe00;
			16'h923a: y = 16'hfe00;
			16'h923b: y = 16'hfe00;
			16'h923c: y = 16'hfe00;
			16'h923d: y = 16'hfe00;
			16'h923e: y = 16'hfe00;
			16'h923f: y = 16'hfe00;
			16'h9240: y = 16'hfe00;
			16'h9241: y = 16'hfe00;
			16'h9242: y = 16'hfe00;
			16'h9243: y = 16'hfe00;
			16'h9244: y = 16'hfe00;
			16'h9245: y = 16'hfe00;
			16'h9246: y = 16'hfe00;
			16'h9247: y = 16'hfe00;
			16'h9248: y = 16'hfe00;
			16'h9249: y = 16'hfe00;
			16'h924a: y = 16'hfe00;
			16'h924b: y = 16'hfe00;
			16'h924c: y = 16'hfe00;
			16'h924d: y = 16'hfe00;
			16'h924e: y = 16'hfe00;
			16'h924f: y = 16'hfe00;
			16'h9250: y = 16'hfe00;
			16'h9251: y = 16'hfe00;
			16'h9252: y = 16'hfe00;
			16'h9253: y = 16'hfe00;
			16'h9254: y = 16'hfe00;
			16'h9255: y = 16'hfe00;
			16'h9256: y = 16'hfe00;
			16'h9257: y = 16'hfe00;
			16'h9258: y = 16'hfe00;
			16'h9259: y = 16'hfe00;
			16'h925a: y = 16'hfe00;
			16'h925b: y = 16'hfe00;
			16'h925c: y = 16'hfe00;
			16'h925d: y = 16'hfe00;
			16'h925e: y = 16'hfe00;
			16'h925f: y = 16'hfe00;
			16'h9260: y = 16'hfe00;
			16'h9261: y = 16'hfe00;
			16'h9262: y = 16'hfe00;
			16'h9263: y = 16'hfe00;
			16'h9264: y = 16'hfe00;
			16'h9265: y = 16'hfe00;
			16'h9266: y = 16'hfe00;
			16'h9267: y = 16'hfe00;
			16'h9268: y = 16'hfe00;
			16'h9269: y = 16'hfe00;
			16'h926a: y = 16'hfe00;
			16'h926b: y = 16'hfe00;
			16'h926c: y = 16'hfe00;
			16'h926d: y = 16'hfe00;
			16'h926e: y = 16'hfe00;
			16'h926f: y = 16'hfe00;
			16'h9270: y = 16'hfe00;
			16'h9271: y = 16'hfe00;
			16'h9272: y = 16'hfe00;
			16'h9273: y = 16'hfe00;
			16'h9274: y = 16'hfe00;
			16'h9275: y = 16'hfe00;
			16'h9276: y = 16'hfe00;
			16'h9277: y = 16'hfe00;
			16'h9278: y = 16'hfe00;
			16'h9279: y = 16'hfe00;
			16'h927a: y = 16'hfe00;
			16'h927b: y = 16'hfe00;
			16'h927c: y = 16'hfe00;
			16'h927d: y = 16'hfe00;
			16'h927e: y = 16'hfe00;
			16'h927f: y = 16'hfe00;
			16'h9280: y = 16'hfe00;
			16'h9281: y = 16'hfe00;
			16'h9282: y = 16'hfe00;
			16'h9283: y = 16'hfe00;
			16'h9284: y = 16'hfe00;
			16'h9285: y = 16'hfe00;
			16'h9286: y = 16'hfe00;
			16'h9287: y = 16'hfe00;
			16'h9288: y = 16'hfe00;
			16'h9289: y = 16'hfe00;
			16'h928a: y = 16'hfe00;
			16'h928b: y = 16'hfe00;
			16'h928c: y = 16'hfe00;
			16'h928d: y = 16'hfe00;
			16'h928e: y = 16'hfe00;
			16'h928f: y = 16'hfe00;
			16'h9290: y = 16'hfe00;
			16'h9291: y = 16'hfe00;
			16'h9292: y = 16'hfe00;
			16'h9293: y = 16'hfe00;
			16'h9294: y = 16'hfe00;
			16'h9295: y = 16'hfe00;
			16'h9296: y = 16'hfe00;
			16'h9297: y = 16'hfe00;
			16'h9298: y = 16'hfe00;
			16'h9299: y = 16'hfe00;
			16'h929a: y = 16'hfe00;
			16'h929b: y = 16'hfe00;
			16'h929c: y = 16'hfe00;
			16'h929d: y = 16'hfe00;
			16'h929e: y = 16'hfe00;
			16'h929f: y = 16'hfe00;
			16'h92a0: y = 16'hfe00;
			16'h92a1: y = 16'hfe00;
			16'h92a2: y = 16'hfe00;
			16'h92a3: y = 16'hfe00;
			16'h92a4: y = 16'hfe00;
			16'h92a5: y = 16'hfe00;
			16'h92a6: y = 16'hfe00;
			16'h92a7: y = 16'hfe00;
			16'h92a8: y = 16'hfe00;
			16'h92a9: y = 16'hfe00;
			16'h92aa: y = 16'hfe00;
			16'h92ab: y = 16'hfe00;
			16'h92ac: y = 16'hfe00;
			16'h92ad: y = 16'hfe00;
			16'h92ae: y = 16'hfe00;
			16'h92af: y = 16'hfe00;
			16'h92b0: y = 16'hfe00;
			16'h92b1: y = 16'hfe00;
			16'h92b2: y = 16'hfe00;
			16'h92b3: y = 16'hfe00;
			16'h92b4: y = 16'hfe00;
			16'h92b5: y = 16'hfe00;
			16'h92b6: y = 16'hfe00;
			16'h92b7: y = 16'hfe00;
			16'h92b8: y = 16'hfe00;
			16'h92b9: y = 16'hfe00;
			16'h92ba: y = 16'hfe00;
			16'h92bb: y = 16'hfe00;
			16'h92bc: y = 16'hfe00;
			16'h92bd: y = 16'hfe00;
			16'h92be: y = 16'hfe00;
			16'h92bf: y = 16'hfe00;
			16'h92c0: y = 16'hfe00;
			16'h92c1: y = 16'hfe00;
			16'h92c2: y = 16'hfe00;
			16'h92c3: y = 16'hfe00;
			16'h92c4: y = 16'hfe00;
			16'h92c5: y = 16'hfe00;
			16'h92c6: y = 16'hfe00;
			16'h92c7: y = 16'hfe00;
			16'h92c8: y = 16'hfe00;
			16'h92c9: y = 16'hfe00;
			16'h92ca: y = 16'hfe00;
			16'h92cb: y = 16'hfe00;
			16'h92cc: y = 16'hfe00;
			16'h92cd: y = 16'hfe00;
			16'h92ce: y = 16'hfe00;
			16'h92cf: y = 16'hfe00;
			16'h92d0: y = 16'hfe00;
			16'h92d1: y = 16'hfe00;
			16'h92d2: y = 16'hfe00;
			16'h92d3: y = 16'hfe00;
			16'h92d4: y = 16'hfe00;
			16'h92d5: y = 16'hfe00;
			16'h92d6: y = 16'hfe00;
			16'h92d7: y = 16'hfe00;
			16'h92d8: y = 16'hfe00;
			16'h92d9: y = 16'hfe00;
			16'h92da: y = 16'hfe00;
			16'h92db: y = 16'hfe00;
			16'h92dc: y = 16'hfe00;
			16'h92dd: y = 16'hfe00;
			16'h92de: y = 16'hfe00;
			16'h92df: y = 16'hfe00;
			16'h92e0: y = 16'hfe00;
			16'h92e1: y = 16'hfe00;
			16'h92e2: y = 16'hfe00;
			16'h92e3: y = 16'hfe00;
			16'h92e4: y = 16'hfe00;
			16'h92e5: y = 16'hfe00;
			16'h92e6: y = 16'hfe00;
			16'h92e7: y = 16'hfe00;
			16'h92e8: y = 16'hfe00;
			16'h92e9: y = 16'hfe00;
			16'h92ea: y = 16'hfe00;
			16'h92eb: y = 16'hfe00;
			16'h92ec: y = 16'hfe00;
			16'h92ed: y = 16'hfe00;
			16'h92ee: y = 16'hfe00;
			16'h92ef: y = 16'hfe00;
			16'h92f0: y = 16'hfe00;
			16'h92f1: y = 16'hfe00;
			16'h92f2: y = 16'hfe00;
			16'h92f3: y = 16'hfe00;
			16'h92f4: y = 16'hfe00;
			16'h92f5: y = 16'hfe00;
			16'h92f6: y = 16'hfe00;
			16'h92f7: y = 16'hfe00;
			16'h92f8: y = 16'hfe00;
			16'h92f9: y = 16'hfe00;
			16'h92fa: y = 16'hfe00;
			16'h92fb: y = 16'hfe00;
			16'h92fc: y = 16'hfe00;
			16'h92fd: y = 16'hfe00;
			16'h92fe: y = 16'hfe00;
			16'h92ff: y = 16'hfe00;
			16'h9300: y = 16'hfe00;
			16'h9301: y = 16'hfe00;
			16'h9302: y = 16'hfe00;
			16'h9303: y = 16'hfe00;
			16'h9304: y = 16'hfe00;
			16'h9305: y = 16'hfe00;
			16'h9306: y = 16'hfe00;
			16'h9307: y = 16'hfe00;
			16'h9308: y = 16'hfe00;
			16'h9309: y = 16'hfe00;
			16'h930a: y = 16'hfe00;
			16'h930b: y = 16'hfe00;
			16'h930c: y = 16'hfe00;
			16'h930d: y = 16'hfe00;
			16'h930e: y = 16'hfe00;
			16'h930f: y = 16'hfe00;
			16'h9310: y = 16'hfe00;
			16'h9311: y = 16'hfe00;
			16'h9312: y = 16'hfe00;
			16'h9313: y = 16'hfe00;
			16'h9314: y = 16'hfe00;
			16'h9315: y = 16'hfe00;
			16'h9316: y = 16'hfe00;
			16'h9317: y = 16'hfe00;
			16'h9318: y = 16'hfe00;
			16'h9319: y = 16'hfe00;
			16'h931a: y = 16'hfe00;
			16'h931b: y = 16'hfe00;
			16'h931c: y = 16'hfe00;
			16'h931d: y = 16'hfe00;
			16'h931e: y = 16'hfe00;
			16'h931f: y = 16'hfe00;
			16'h9320: y = 16'hfe00;
			16'h9321: y = 16'hfe00;
			16'h9322: y = 16'hfe00;
			16'h9323: y = 16'hfe00;
			16'h9324: y = 16'hfe00;
			16'h9325: y = 16'hfe00;
			16'h9326: y = 16'hfe00;
			16'h9327: y = 16'hfe00;
			16'h9328: y = 16'hfe00;
			16'h9329: y = 16'hfe00;
			16'h932a: y = 16'hfe00;
			16'h932b: y = 16'hfe00;
			16'h932c: y = 16'hfe00;
			16'h932d: y = 16'hfe00;
			16'h932e: y = 16'hfe00;
			16'h932f: y = 16'hfe00;
			16'h9330: y = 16'hfe00;
			16'h9331: y = 16'hfe00;
			16'h9332: y = 16'hfe00;
			16'h9333: y = 16'hfe00;
			16'h9334: y = 16'hfe00;
			16'h9335: y = 16'hfe00;
			16'h9336: y = 16'hfe00;
			16'h9337: y = 16'hfe00;
			16'h9338: y = 16'hfe00;
			16'h9339: y = 16'hfe00;
			16'h933a: y = 16'hfe00;
			16'h933b: y = 16'hfe00;
			16'h933c: y = 16'hfe00;
			16'h933d: y = 16'hfe00;
			16'h933e: y = 16'hfe00;
			16'h933f: y = 16'hfe00;
			16'h9340: y = 16'hfe00;
			16'h9341: y = 16'hfe00;
			16'h9342: y = 16'hfe00;
			16'h9343: y = 16'hfe00;
			16'h9344: y = 16'hfe00;
			16'h9345: y = 16'hfe00;
			16'h9346: y = 16'hfe00;
			16'h9347: y = 16'hfe00;
			16'h9348: y = 16'hfe00;
			16'h9349: y = 16'hfe00;
			16'h934a: y = 16'hfe00;
			16'h934b: y = 16'hfe00;
			16'h934c: y = 16'hfe00;
			16'h934d: y = 16'hfe00;
			16'h934e: y = 16'hfe00;
			16'h934f: y = 16'hfe00;
			16'h9350: y = 16'hfe00;
			16'h9351: y = 16'hfe00;
			16'h9352: y = 16'hfe00;
			16'h9353: y = 16'hfe00;
			16'h9354: y = 16'hfe00;
			16'h9355: y = 16'hfe00;
			16'h9356: y = 16'hfe00;
			16'h9357: y = 16'hfe00;
			16'h9358: y = 16'hfe00;
			16'h9359: y = 16'hfe00;
			16'h935a: y = 16'hfe00;
			16'h935b: y = 16'hfe00;
			16'h935c: y = 16'hfe00;
			16'h935d: y = 16'hfe00;
			16'h935e: y = 16'hfe00;
			16'h935f: y = 16'hfe00;
			16'h9360: y = 16'hfe00;
			16'h9361: y = 16'hfe00;
			16'h9362: y = 16'hfe00;
			16'h9363: y = 16'hfe00;
			16'h9364: y = 16'hfe00;
			16'h9365: y = 16'hfe00;
			16'h9366: y = 16'hfe00;
			16'h9367: y = 16'hfe00;
			16'h9368: y = 16'hfe00;
			16'h9369: y = 16'hfe00;
			16'h936a: y = 16'hfe00;
			16'h936b: y = 16'hfe00;
			16'h936c: y = 16'hfe00;
			16'h936d: y = 16'hfe00;
			16'h936e: y = 16'hfe00;
			16'h936f: y = 16'hfe00;
			16'h9370: y = 16'hfe00;
			16'h9371: y = 16'hfe00;
			16'h9372: y = 16'hfe00;
			16'h9373: y = 16'hfe00;
			16'h9374: y = 16'hfe00;
			16'h9375: y = 16'hfe00;
			16'h9376: y = 16'hfe00;
			16'h9377: y = 16'hfe00;
			16'h9378: y = 16'hfe00;
			16'h9379: y = 16'hfe00;
			16'h937a: y = 16'hfe00;
			16'h937b: y = 16'hfe00;
			16'h937c: y = 16'hfe00;
			16'h937d: y = 16'hfe00;
			16'h937e: y = 16'hfe00;
			16'h937f: y = 16'hfe00;
			16'h9380: y = 16'hfe00;
			16'h9381: y = 16'hfe00;
			16'h9382: y = 16'hfe00;
			16'h9383: y = 16'hfe00;
			16'h9384: y = 16'hfe00;
			16'h9385: y = 16'hfe00;
			16'h9386: y = 16'hfe00;
			16'h9387: y = 16'hfe00;
			16'h9388: y = 16'hfe00;
			16'h9389: y = 16'hfe00;
			16'h938a: y = 16'hfe00;
			16'h938b: y = 16'hfe00;
			16'h938c: y = 16'hfe00;
			16'h938d: y = 16'hfe00;
			16'h938e: y = 16'hfe00;
			16'h938f: y = 16'hfe00;
			16'h9390: y = 16'hfe00;
			16'h9391: y = 16'hfe00;
			16'h9392: y = 16'hfe00;
			16'h9393: y = 16'hfe00;
			16'h9394: y = 16'hfe00;
			16'h9395: y = 16'hfe00;
			16'h9396: y = 16'hfe00;
			16'h9397: y = 16'hfe00;
			16'h9398: y = 16'hfe00;
			16'h9399: y = 16'hfe00;
			16'h939a: y = 16'hfe00;
			16'h939b: y = 16'hfe00;
			16'h939c: y = 16'hfe00;
			16'h939d: y = 16'hfe00;
			16'h939e: y = 16'hfe00;
			16'h939f: y = 16'hfe00;
			16'h93a0: y = 16'hfe00;
			16'h93a1: y = 16'hfe00;
			16'h93a2: y = 16'hfe00;
			16'h93a3: y = 16'hfe00;
			16'h93a4: y = 16'hfe00;
			16'h93a5: y = 16'hfe00;
			16'h93a6: y = 16'hfe00;
			16'h93a7: y = 16'hfe00;
			16'h93a8: y = 16'hfe00;
			16'h93a9: y = 16'hfe00;
			16'h93aa: y = 16'hfe00;
			16'h93ab: y = 16'hfe00;
			16'h93ac: y = 16'hfe00;
			16'h93ad: y = 16'hfe00;
			16'h93ae: y = 16'hfe00;
			16'h93af: y = 16'hfe00;
			16'h93b0: y = 16'hfe00;
			16'h93b1: y = 16'hfe00;
			16'h93b2: y = 16'hfe00;
			16'h93b3: y = 16'hfe00;
			16'h93b4: y = 16'hfe00;
			16'h93b5: y = 16'hfe00;
			16'h93b6: y = 16'hfe00;
			16'h93b7: y = 16'hfe00;
			16'h93b8: y = 16'hfe00;
			16'h93b9: y = 16'hfe00;
			16'h93ba: y = 16'hfe00;
			16'h93bb: y = 16'hfe00;
			16'h93bc: y = 16'hfe00;
			16'h93bd: y = 16'hfe00;
			16'h93be: y = 16'hfe00;
			16'h93bf: y = 16'hfe00;
			16'h93c0: y = 16'hfe00;
			16'h93c1: y = 16'hfe00;
			16'h93c2: y = 16'hfe00;
			16'h93c3: y = 16'hfe00;
			16'h93c4: y = 16'hfe00;
			16'h93c5: y = 16'hfe00;
			16'h93c6: y = 16'hfe00;
			16'h93c7: y = 16'hfe00;
			16'h93c8: y = 16'hfe00;
			16'h93c9: y = 16'hfe00;
			16'h93ca: y = 16'hfe00;
			16'h93cb: y = 16'hfe00;
			16'h93cc: y = 16'hfe00;
			16'h93cd: y = 16'hfe00;
			16'h93ce: y = 16'hfe00;
			16'h93cf: y = 16'hfe00;
			16'h93d0: y = 16'hfe00;
			16'h93d1: y = 16'hfe00;
			16'h93d2: y = 16'hfe00;
			16'h93d3: y = 16'hfe00;
			16'h93d4: y = 16'hfe00;
			16'h93d5: y = 16'hfe00;
			16'h93d6: y = 16'hfe00;
			16'h93d7: y = 16'hfe00;
			16'h93d8: y = 16'hfe00;
			16'h93d9: y = 16'hfe00;
			16'h93da: y = 16'hfe00;
			16'h93db: y = 16'hfe00;
			16'h93dc: y = 16'hfe00;
			16'h93dd: y = 16'hfe00;
			16'h93de: y = 16'hfe00;
			16'h93df: y = 16'hfe00;
			16'h93e0: y = 16'hfe00;
			16'h93e1: y = 16'hfe00;
			16'h93e2: y = 16'hfe00;
			16'h93e3: y = 16'hfe00;
			16'h93e4: y = 16'hfe00;
			16'h93e5: y = 16'hfe00;
			16'h93e6: y = 16'hfe00;
			16'h93e7: y = 16'hfe00;
			16'h93e8: y = 16'hfe00;
			16'h93e9: y = 16'hfe00;
			16'h93ea: y = 16'hfe00;
			16'h93eb: y = 16'hfe00;
			16'h93ec: y = 16'hfe00;
			16'h93ed: y = 16'hfe00;
			16'h93ee: y = 16'hfe00;
			16'h93ef: y = 16'hfe00;
			16'h93f0: y = 16'hfe00;
			16'h93f1: y = 16'hfe00;
			16'h93f2: y = 16'hfe00;
			16'h93f3: y = 16'hfe00;
			16'h93f4: y = 16'hfe00;
			16'h93f5: y = 16'hfe00;
			16'h93f6: y = 16'hfe00;
			16'h93f7: y = 16'hfe00;
			16'h93f8: y = 16'hfe00;
			16'h93f9: y = 16'hfe00;
			16'h93fa: y = 16'hfe00;
			16'h93fb: y = 16'hfe00;
			16'h93fc: y = 16'hfe00;
			16'h93fd: y = 16'hfe00;
			16'h93fe: y = 16'hfe00;
			16'h93ff: y = 16'hfe00;
			16'h9400: y = 16'hfe00;
			16'h9401: y = 16'hfe00;
			16'h9402: y = 16'hfe00;
			16'h9403: y = 16'hfe00;
			16'h9404: y = 16'hfe00;
			16'h9405: y = 16'hfe00;
			16'h9406: y = 16'hfe00;
			16'h9407: y = 16'hfe00;
			16'h9408: y = 16'hfe00;
			16'h9409: y = 16'hfe00;
			16'h940a: y = 16'hfe00;
			16'h940b: y = 16'hfe00;
			16'h940c: y = 16'hfe00;
			16'h940d: y = 16'hfe00;
			16'h940e: y = 16'hfe00;
			16'h940f: y = 16'hfe00;
			16'h9410: y = 16'hfe00;
			16'h9411: y = 16'hfe00;
			16'h9412: y = 16'hfe00;
			16'h9413: y = 16'hfe00;
			16'h9414: y = 16'hfe00;
			16'h9415: y = 16'hfe00;
			16'h9416: y = 16'hfe00;
			16'h9417: y = 16'hfe00;
			16'h9418: y = 16'hfe00;
			16'h9419: y = 16'hfe00;
			16'h941a: y = 16'hfe00;
			16'h941b: y = 16'hfe00;
			16'h941c: y = 16'hfe00;
			16'h941d: y = 16'hfe00;
			16'h941e: y = 16'hfe00;
			16'h941f: y = 16'hfe00;
			16'h9420: y = 16'hfe00;
			16'h9421: y = 16'hfe00;
			16'h9422: y = 16'hfe00;
			16'h9423: y = 16'hfe00;
			16'h9424: y = 16'hfe00;
			16'h9425: y = 16'hfe00;
			16'h9426: y = 16'hfe00;
			16'h9427: y = 16'hfe00;
			16'h9428: y = 16'hfe00;
			16'h9429: y = 16'hfe00;
			16'h942a: y = 16'hfe00;
			16'h942b: y = 16'hfe00;
			16'h942c: y = 16'hfe00;
			16'h942d: y = 16'hfe00;
			16'h942e: y = 16'hfe00;
			16'h942f: y = 16'hfe00;
			16'h9430: y = 16'hfe00;
			16'h9431: y = 16'hfe00;
			16'h9432: y = 16'hfe00;
			16'h9433: y = 16'hfe00;
			16'h9434: y = 16'hfe00;
			16'h9435: y = 16'hfe00;
			16'h9436: y = 16'hfe00;
			16'h9437: y = 16'hfe00;
			16'h9438: y = 16'hfe00;
			16'h9439: y = 16'hfe00;
			16'h943a: y = 16'hfe00;
			16'h943b: y = 16'hfe00;
			16'h943c: y = 16'hfe00;
			16'h943d: y = 16'hfe00;
			16'h943e: y = 16'hfe00;
			16'h943f: y = 16'hfe00;
			16'h9440: y = 16'hfe00;
			16'h9441: y = 16'hfe00;
			16'h9442: y = 16'hfe00;
			16'h9443: y = 16'hfe00;
			16'h9444: y = 16'hfe00;
			16'h9445: y = 16'hfe00;
			16'h9446: y = 16'hfe00;
			16'h9447: y = 16'hfe00;
			16'h9448: y = 16'hfe00;
			16'h9449: y = 16'hfe00;
			16'h944a: y = 16'hfe00;
			16'h944b: y = 16'hfe00;
			16'h944c: y = 16'hfe00;
			16'h944d: y = 16'hfe00;
			16'h944e: y = 16'hfe00;
			16'h944f: y = 16'hfe00;
			16'h9450: y = 16'hfe00;
			16'h9451: y = 16'hfe00;
			16'h9452: y = 16'hfe00;
			16'h9453: y = 16'hfe00;
			16'h9454: y = 16'hfe00;
			16'h9455: y = 16'hfe00;
			16'h9456: y = 16'hfe00;
			16'h9457: y = 16'hfe00;
			16'h9458: y = 16'hfe00;
			16'h9459: y = 16'hfe00;
			16'h945a: y = 16'hfe00;
			16'h945b: y = 16'hfe00;
			16'h945c: y = 16'hfe00;
			16'h945d: y = 16'hfe00;
			16'h945e: y = 16'hfe00;
			16'h945f: y = 16'hfe00;
			16'h9460: y = 16'hfe00;
			16'h9461: y = 16'hfe00;
			16'h9462: y = 16'hfe00;
			16'h9463: y = 16'hfe00;
			16'h9464: y = 16'hfe00;
			16'h9465: y = 16'hfe00;
			16'h9466: y = 16'hfe00;
			16'h9467: y = 16'hfe00;
			16'h9468: y = 16'hfe00;
			16'h9469: y = 16'hfe00;
			16'h946a: y = 16'hfe00;
			16'h946b: y = 16'hfe00;
			16'h946c: y = 16'hfe00;
			16'h946d: y = 16'hfe00;
			16'h946e: y = 16'hfe00;
			16'h946f: y = 16'hfe00;
			16'h9470: y = 16'hfe00;
			16'h9471: y = 16'hfe00;
			16'h9472: y = 16'hfe00;
			16'h9473: y = 16'hfe00;
			16'h9474: y = 16'hfe00;
			16'h9475: y = 16'hfe00;
			16'h9476: y = 16'hfe00;
			16'h9477: y = 16'hfe00;
			16'h9478: y = 16'hfe00;
			16'h9479: y = 16'hfe00;
			16'h947a: y = 16'hfe00;
			16'h947b: y = 16'hfe00;
			16'h947c: y = 16'hfe00;
			16'h947d: y = 16'hfe00;
			16'h947e: y = 16'hfe00;
			16'h947f: y = 16'hfe00;
			16'h9480: y = 16'hfe00;
			16'h9481: y = 16'hfe00;
			16'h9482: y = 16'hfe00;
			16'h9483: y = 16'hfe00;
			16'h9484: y = 16'hfe00;
			16'h9485: y = 16'hfe00;
			16'h9486: y = 16'hfe00;
			16'h9487: y = 16'hfe00;
			16'h9488: y = 16'hfe00;
			16'h9489: y = 16'hfe00;
			16'h948a: y = 16'hfe00;
			16'h948b: y = 16'hfe00;
			16'h948c: y = 16'hfe00;
			16'h948d: y = 16'hfe00;
			16'h948e: y = 16'hfe00;
			16'h948f: y = 16'hfe00;
			16'h9490: y = 16'hfe00;
			16'h9491: y = 16'hfe00;
			16'h9492: y = 16'hfe00;
			16'h9493: y = 16'hfe00;
			16'h9494: y = 16'hfe00;
			16'h9495: y = 16'hfe00;
			16'h9496: y = 16'hfe00;
			16'h9497: y = 16'hfe00;
			16'h9498: y = 16'hfe00;
			16'h9499: y = 16'hfe00;
			16'h949a: y = 16'hfe00;
			16'h949b: y = 16'hfe00;
			16'h949c: y = 16'hfe00;
			16'h949d: y = 16'hfe00;
			16'h949e: y = 16'hfe00;
			16'h949f: y = 16'hfe00;
			16'h94a0: y = 16'hfe00;
			16'h94a1: y = 16'hfe00;
			16'h94a2: y = 16'hfe00;
			16'h94a3: y = 16'hfe00;
			16'h94a4: y = 16'hfe00;
			16'h94a5: y = 16'hfe00;
			16'h94a6: y = 16'hfe00;
			16'h94a7: y = 16'hfe00;
			16'h94a8: y = 16'hfe00;
			16'h94a9: y = 16'hfe00;
			16'h94aa: y = 16'hfe00;
			16'h94ab: y = 16'hfe00;
			16'h94ac: y = 16'hfe00;
			16'h94ad: y = 16'hfe00;
			16'h94ae: y = 16'hfe00;
			16'h94af: y = 16'hfe00;
			16'h94b0: y = 16'hfe00;
			16'h94b1: y = 16'hfe00;
			16'h94b2: y = 16'hfe00;
			16'h94b3: y = 16'hfe00;
			16'h94b4: y = 16'hfe00;
			16'h94b5: y = 16'hfe00;
			16'h94b6: y = 16'hfe00;
			16'h94b7: y = 16'hfe00;
			16'h94b8: y = 16'hfe00;
			16'h94b9: y = 16'hfe00;
			16'h94ba: y = 16'hfe00;
			16'h94bb: y = 16'hfe00;
			16'h94bc: y = 16'hfe00;
			16'h94bd: y = 16'hfe00;
			16'h94be: y = 16'hfe00;
			16'h94bf: y = 16'hfe00;
			16'h94c0: y = 16'hfe00;
			16'h94c1: y = 16'hfe00;
			16'h94c2: y = 16'hfe00;
			16'h94c3: y = 16'hfe00;
			16'h94c4: y = 16'hfe00;
			16'h94c5: y = 16'hfe00;
			16'h94c6: y = 16'hfe00;
			16'h94c7: y = 16'hfe00;
			16'h94c8: y = 16'hfe00;
			16'h94c9: y = 16'hfe00;
			16'h94ca: y = 16'hfe00;
			16'h94cb: y = 16'hfe00;
			16'h94cc: y = 16'hfe00;
			16'h94cd: y = 16'hfe00;
			16'h94ce: y = 16'hfe00;
			16'h94cf: y = 16'hfe00;
			16'h94d0: y = 16'hfe00;
			16'h94d1: y = 16'hfe00;
			16'h94d2: y = 16'hfe00;
			16'h94d3: y = 16'hfe00;
			16'h94d4: y = 16'hfe00;
			16'h94d5: y = 16'hfe00;
			16'h94d6: y = 16'hfe00;
			16'h94d7: y = 16'hfe00;
			16'h94d8: y = 16'hfe00;
			16'h94d9: y = 16'hfe00;
			16'h94da: y = 16'hfe00;
			16'h94db: y = 16'hfe00;
			16'h94dc: y = 16'hfe00;
			16'h94dd: y = 16'hfe00;
			16'h94de: y = 16'hfe00;
			16'h94df: y = 16'hfe00;
			16'h94e0: y = 16'hfe00;
			16'h94e1: y = 16'hfe00;
			16'h94e2: y = 16'hfe00;
			16'h94e3: y = 16'hfe00;
			16'h94e4: y = 16'hfe00;
			16'h94e5: y = 16'hfe00;
			16'h94e6: y = 16'hfe00;
			16'h94e7: y = 16'hfe00;
			16'h94e8: y = 16'hfe00;
			16'h94e9: y = 16'hfe00;
			16'h94ea: y = 16'hfe00;
			16'h94eb: y = 16'hfe00;
			16'h94ec: y = 16'hfe00;
			16'h94ed: y = 16'hfe00;
			16'h94ee: y = 16'hfe00;
			16'h94ef: y = 16'hfe00;
			16'h94f0: y = 16'hfe00;
			16'h94f1: y = 16'hfe00;
			16'h94f2: y = 16'hfe00;
			16'h94f3: y = 16'hfe00;
			16'h94f4: y = 16'hfe00;
			16'h94f5: y = 16'hfe00;
			16'h94f6: y = 16'hfe00;
			16'h94f7: y = 16'hfe00;
			16'h94f8: y = 16'hfe00;
			16'h94f9: y = 16'hfe00;
			16'h94fa: y = 16'hfe00;
			16'h94fb: y = 16'hfe00;
			16'h94fc: y = 16'hfe00;
			16'h94fd: y = 16'hfe00;
			16'h94fe: y = 16'hfe00;
			16'h94ff: y = 16'hfe00;
			16'h9500: y = 16'hfe00;
			16'h9501: y = 16'hfe00;
			16'h9502: y = 16'hfe00;
			16'h9503: y = 16'hfe00;
			16'h9504: y = 16'hfe00;
			16'h9505: y = 16'hfe00;
			16'h9506: y = 16'hfe00;
			16'h9507: y = 16'hfe00;
			16'h9508: y = 16'hfe00;
			16'h9509: y = 16'hfe00;
			16'h950a: y = 16'hfe00;
			16'h950b: y = 16'hfe00;
			16'h950c: y = 16'hfe00;
			16'h950d: y = 16'hfe00;
			16'h950e: y = 16'hfe00;
			16'h950f: y = 16'hfe00;
			16'h9510: y = 16'hfe00;
			16'h9511: y = 16'hfe00;
			16'h9512: y = 16'hfe00;
			16'h9513: y = 16'hfe00;
			16'h9514: y = 16'hfe00;
			16'h9515: y = 16'hfe00;
			16'h9516: y = 16'hfe00;
			16'h9517: y = 16'hfe00;
			16'h9518: y = 16'hfe00;
			16'h9519: y = 16'hfe00;
			16'h951a: y = 16'hfe00;
			16'h951b: y = 16'hfe00;
			16'h951c: y = 16'hfe00;
			16'h951d: y = 16'hfe00;
			16'h951e: y = 16'hfe00;
			16'h951f: y = 16'hfe00;
			16'h9520: y = 16'hfe00;
			16'h9521: y = 16'hfe00;
			16'h9522: y = 16'hfe00;
			16'h9523: y = 16'hfe00;
			16'h9524: y = 16'hfe00;
			16'h9525: y = 16'hfe00;
			16'h9526: y = 16'hfe00;
			16'h9527: y = 16'hfe00;
			16'h9528: y = 16'hfe00;
			16'h9529: y = 16'hfe00;
			16'h952a: y = 16'hfe00;
			16'h952b: y = 16'hfe00;
			16'h952c: y = 16'hfe00;
			16'h952d: y = 16'hfe00;
			16'h952e: y = 16'hfe00;
			16'h952f: y = 16'hfe00;
			16'h9530: y = 16'hfe00;
			16'h9531: y = 16'hfe00;
			16'h9532: y = 16'hfe00;
			16'h9533: y = 16'hfe00;
			16'h9534: y = 16'hfe00;
			16'h9535: y = 16'hfe00;
			16'h9536: y = 16'hfe00;
			16'h9537: y = 16'hfe00;
			16'h9538: y = 16'hfe00;
			16'h9539: y = 16'hfe00;
			16'h953a: y = 16'hfe00;
			16'h953b: y = 16'hfe00;
			16'h953c: y = 16'hfe00;
			16'h953d: y = 16'hfe00;
			16'h953e: y = 16'hfe00;
			16'h953f: y = 16'hfe00;
			16'h9540: y = 16'hfe00;
			16'h9541: y = 16'hfe00;
			16'h9542: y = 16'hfe00;
			16'h9543: y = 16'hfe00;
			16'h9544: y = 16'hfe00;
			16'h9545: y = 16'hfe00;
			16'h9546: y = 16'hfe00;
			16'h9547: y = 16'hfe00;
			16'h9548: y = 16'hfe00;
			16'h9549: y = 16'hfe00;
			16'h954a: y = 16'hfe00;
			16'h954b: y = 16'hfe00;
			16'h954c: y = 16'hfe00;
			16'h954d: y = 16'hfe00;
			16'h954e: y = 16'hfe00;
			16'h954f: y = 16'hfe00;
			16'h9550: y = 16'hfe00;
			16'h9551: y = 16'hfe00;
			16'h9552: y = 16'hfe00;
			16'h9553: y = 16'hfe00;
			16'h9554: y = 16'hfe00;
			16'h9555: y = 16'hfe00;
			16'h9556: y = 16'hfe00;
			16'h9557: y = 16'hfe00;
			16'h9558: y = 16'hfe00;
			16'h9559: y = 16'hfe00;
			16'h955a: y = 16'hfe00;
			16'h955b: y = 16'hfe00;
			16'h955c: y = 16'hfe00;
			16'h955d: y = 16'hfe00;
			16'h955e: y = 16'hfe00;
			16'h955f: y = 16'hfe00;
			16'h9560: y = 16'hfe00;
			16'h9561: y = 16'hfe00;
			16'h9562: y = 16'hfe00;
			16'h9563: y = 16'hfe00;
			16'h9564: y = 16'hfe00;
			16'h9565: y = 16'hfe00;
			16'h9566: y = 16'hfe00;
			16'h9567: y = 16'hfe00;
			16'h9568: y = 16'hfe00;
			16'h9569: y = 16'hfe00;
			16'h956a: y = 16'hfe00;
			16'h956b: y = 16'hfe00;
			16'h956c: y = 16'hfe00;
			16'h956d: y = 16'hfe00;
			16'h956e: y = 16'hfe00;
			16'h956f: y = 16'hfe00;
			16'h9570: y = 16'hfe00;
			16'h9571: y = 16'hfe00;
			16'h9572: y = 16'hfe00;
			16'h9573: y = 16'hfe00;
			16'h9574: y = 16'hfe00;
			16'h9575: y = 16'hfe00;
			16'h9576: y = 16'hfe00;
			16'h9577: y = 16'hfe00;
			16'h9578: y = 16'hfe00;
			16'h9579: y = 16'hfe00;
			16'h957a: y = 16'hfe00;
			16'h957b: y = 16'hfe00;
			16'h957c: y = 16'hfe00;
			16'h957d: y = 16'hfe00;
			16'h957e: y = 16'hfe00;
			16'h957f: y = 16'hfe00;
			16'h9580: y = 16'hfe00;
			16'h9581: y = 16'hfe00;
			16'h9582: y = 16'hfe00;
			16'h9583: y = 16'hfe00;
			16'h9584: y = 16'hfe00;
			16'h9585: y = 16'hfe00;
			16'h9586: y = 16'hfe00;
			16'h9587: y = 16'hfe00;
			16'h9588: y = 16'hfe00;
			16'h9589: y = 16'hfe00;
			16'h958a: y = 16'hfe00;
			16'h958b: y = 16'hfe00;
			16'h958c: y = 16'hfe00;
			16'h958d: y = 16'hfe00;
			16'h958e: y = 16'hfe00;
			16'h958f: y = 16'hfe00;
			16'h9590: y = 16'hfe00;
			16'h9591: y = 16'hfe00;
			16'h9592: y = 16'hfe00;
			16'h9593: y = 16'hfe00;
			16'h9594: y = 16'hfe00;
			16'h9595: y = 16'hfe00;
			16'h9596: y = 16'hfe00;
			16'h9597: y = 16'hfe00;
			16'h9598: y = 16'hfe00;
			16'h9599: y = 16'hfe00;
			16'h959a: y = 16'hfe00;
			16'h959b: y = 16'hfe00;
			16'h959c: y = 16'hfe00;
			16'h959d: y = 16'hfe00;
			16'h959e: y = 16'hfe00;
			16'h959f: y = 16'hfe00;
			16'h95a0: y = 16'hfe00;
			16'h95a1: y = 16'hfe00;
			16'h95a2: y = 16'hfe00;
			16'h95a3: y = 16'hfe00;
			16'h95a4: y = 16'hfe00;
			16'h95a5: y = 16'hfe00;
			16'h95a6: y = 16'hfe00;
			16'h95a7: y = 16'hfe00;
			16'h95a8: y = 16'hfe00;
			16'h95a9: y = 16'hfe00;
			16'h95aa: y = 16'hfe00;
			16'h95ab: y = 16'hfe00;
			16'h95ac: y = 16'hfe00;
			16'h95ad: y = 16'hfe00;
			16'h95ae: y = 16'hfe00;
			16'h95af: y = 16'hfe00;
			16'h95b0: y = 16'hfe00;
			16'h95b1: y = 16'hfe00;
			16'h95b2: y = 16'hfe00;
			16'h95b3: y = 16'hfe00;
			16'h95b4: y = 16'hfe00;
			16'h95b5: y = 16'hfe00;
			16'h95b6: y = 16'hfe00;
			16'h95b7: y = 16'hfe00;
			16'h95b8: y = 16'hfe00;
			16'h95b9: y = 16'hfe00;
			16'h95ba: y = 16'hfe00;
			16'h95bb: y = 16'hfe00;
			16'h95bc: y = 16'hfe00;
			16'h95bd: y = 16'hfe00;
			16'h95be: y = 16'hfe00;
			16'h95bf: y = 16'hfe00;
			16'h95c0: y = 16'hfe00;
			16'h95c1: y = 16'hfe00;
			16'h95c2: y = 16'hfe00;
			16'h95c3: y = 16'hfe00;
			16'h95c4: y = 16'hfe00;
			16'h95c5: y = 16'hfe00;
			16'h95c6: y = 16'hfe00;
			16'h95c7: y = 16'hfe00;
			16'h95c8: y = 16'hfe00;
			16'h95c9: y = 16'hfe00;
			16'h95ca: y = 16'hfe00;
			16'h95cb: y = 16'hfe00;
			16'h95cc: y = 16'hfe00;
			16'h95cd: y = 16'hfe00;
			16'h95ce: y = 16'hfe00;
			16'h95cf: y = 16'hfe00;
			16'h95d0: y = 16'hfe00;
			16'h95d1: y = 16'hfe00;
			16'h95d2: y = 16'hfe00;
			16'h95d3: y = 16'hfe00;
			16'h95d4: y = 16'hfe00;
			16'h95d5: y = 16'hfe00;
			16'h95d6: y = 16'hfe00;
			16'h95d7: y = 16'hfe00;
			16'h95d8: y = 16'hfe00;
			16'h95d9: y = 16'hfe00;
			16'h95da: y = 16'hfe00;
			16'h95db: y = 16'hfe00;
			16'h95dc: y = 16'hfe00;
			16'h95dd: y = 16'hfe00;
			16'h95de: y = 16'hfe00;
			16'h95df: y = 16'hfe00;
			16'h95e0: y = 16'hfe00;
			16'h95e1: y = 16'hfe00;
			16'h95e2: y = 16'hfe00;
			16'h95e3: y = 16'hfe00;
			16'h95e4: y = 16'hfe00;
			16'h95e5: y = 16'hfe00;
			16'h95e6: y = 16'hfe00;
			16'h95e7: y = 16'hfe00;
			16'h95e8: y = 16'hfe00;
			16'h95e9: y = 16'hfe00;
			16'h95ea: y = 16'hfe00;
			16'h95eb: y = 16'hfe00;
			16'h95ec: y = 16'hfe00;
			16'h95ed: y = 16'hfe00;
			16'h95ee: y = 16'hfe00;
			16'h95ef: y = 16'hfe00;
			16'h95f0: y = 16'hfe00;
			16'h95f1: y = 16'hfe00;
			16'h95f2: y = 16'hfe00;
			16'h95f3: y = 16'hfe00;
			16'h95f4: y = 16'hfe00;
			16'h95f5: y = 16'hfe00;
			16'h95f6: y = 16'hfe00;
			16'h95f7: y = 16'hfe00;
			16'h95f8: y = 16'hfe00;
			16'h95f9: y = 16'hfe00;
			16'h95fa: y = 16'hfe00;
			16'h95fb: y = 16'hfe00;
			16'h95fc: y = 16'hfe00;
			16'h95fd: y = 16'hfe00;
			16'h95fe: y = 16'hfe00;
			16'h95ff: y = 16'hfe00;
			16'h9600: y = 16'hfe00;
			16'h9601: y = 16'hfe00;
			16'h9602: y = 16'hfe00;
			16'h9603: y = 16'hfe00;
			16'h9604: y = 16'hfe00;
			16'h9605: y = 16'hfe00;
			16'h9606: y = 16'hfe00;
			16'h9607: y = 16'hfe00;
			16'h9608: y = 16'hfe00;
			16'h9609: y = 16'hfe00;
			16'h960a: y = 16'hfe00;
			16'h960b: y = 16'hfe00;
			16'h960c: y = 16'hfe00;
			16'h960d: y = 16'hfe00;
			16'h960e: y = 16'hfe00;
			16'h960f: y = 16'hfe00;
			16'h9610: y = 16'hfe00;
			16'h9611: y = 16'hfe00;
			16'h9612: y = 16'hfe00;
			16'h9613: y = 16'hfe00;
			16'h9614: y = 16'hfe00;
			16'h9615: y = 16'hfe00;
			16'h9616: y = 16'hfe00;
			16'h9617: y = 16'hfe00;
			16'h9618: y = 16'hfe00;
			16'h9619: y = 16'hfe00;
			16'h961a: y = 16'hfe00;
			16'h961b: y = 16'hfe00;
			16'h961c: y = 16'hfe00;
			16'h961d: y = 16'hfe00;
			16'h961e: y = 16'hfe00;
			16'h961f: y = 16'hfe00;
			16'h9620: y = 16'hfe00;
			16'h9621: y = 16'hfe00;
			16'h9622: y = 16'hfe00;
			16'h9623: y = 16'hfe00;
			16'h9624: y = 16'hfe00;
			16'h9625: y = 16'hfe00;
			16'h9626: y = 16'hfe00;
			16'h9627: y = 16'hfe00;
			16'h9628: y = 16'hfe00;
			16'h9629: y = 16'hfe00;
			16'h962a: y = 16'hfe00;
			16'h962b: y = 16'hfe00;
			16'h962c: y = 16'hfe00;
			16'h962d: y = 16'hfe00;
			16'h962e: y = 16'hfe00;
			16'h962f: y = 16'hfe00;
			16'h9630: y = 16'hfe00;
			16'h9631: y = 16'hfe00;
			16'h9632: y = 16'hfe00;
			16'h9633: y = 16'hfe00;
			16'h9634: y = 16'hfe00;
			16'h9635: y = 16'hfe00;
			16'h9636: y = 16'hfe00;
			16'h9637: y = 16'hfe00;
			16'h9638: y = 16'hfe00;
			16'h9639: y = 16'hfe00;
			16'h963a: y = 16'hfe00;
			16'h963b: y = 16'hfe00;
			16'h963c: y = 16'hfe00;
			16'h963d: y = 16'hfe00;
			16'h963e: y = 16'hfe00;
			16'h963f: y = 16'hfe00;
			16'h9640: y = 16'hfe00;
			16'h9641: y = 16'hfe00;
			16'h9642: y = 16'hfe00;
			16'h9643: y = 16'hfe00;
			16'h9644: y = 16'hfe00;
			16'h9645: y = 16'hfe00;
			16'h9646: y = 16'hfe00;
			16'h9647: y = 16'hfe00;
			16'h9648: y = 16'hfe00;
			16'h9649: y = 16'hfe00;
			16'h964a: y = 16'hfe00;
			16'h964b: y = 16'hfe00;
			16'h964c: y = 16'hfe00;
			16'h964d: y = 16'hfe00;
			16'h964e: y = 16'hfe00;
			16'h964f: y = 16'hfe00;
			16'h9650: y = 16'hfe00;
			16'h9651: y = 16'hfe00;
			16'h9652: y = 16'hfe00;
			16'h9653: y = 16'hfe00;
			16'h9654: y = 16'hfe00;
			16'h9655: y = 16'hfe00;
			16'h9656: y = 16'hfe00;
			16'h9657: y = 16'hfe00;
			16'h9658: y = 16'hfe00;
			16'h9659: y = 16'hfe00;
			16'h965a: y = 16'hfe00;
			16'h965b: y = 16'hfe00;
			16'h965c: y = 16'hfe00;
			16'h965d: y = 16'hfe00;
			16'h965e: y = 16'hfe00;
			16'h965f: y = 16'hfe00;
			16'h9660: y = 16'hfe00;
			16'h9661: y = 16'hfe00;
			16'h9662: y = 16'hfe00;
			16'h9663: y = 16'hfe00;
			16'h9664: y = 16'hfe00;
			16'h9665: y = 16'hfe00;
			16'h9666: y = 16'hfe00;
			16'h9667: y = 16'hfe00;
			16'h9668: y = 16'hfe00;
			16'h9669: y = 16'hfe00;
			16'h966a: y = 16'hfe00;
			16'h966b: y = 16'hfe00;
			16'h966c: y = 16'hfe00;
			16'h966d: y = 16'hfe00;
			16'h966e: y = 16'hfe00;
			16'h966f: y = 16'hfe00;
			16'h9670: y = 16'hfe00;
			16'h9671: y = 16'hfe00;
			16'h9672: y = 16'hfe00;
			16'h9673: y = 16'hfe00;
			16'h9674: y = 16'hfe00;
			16'h9675: y = 16'hfe00;
			16'h9676: y = 16'hfe00;
			16'h9677: y = 16'hfe00;
			16'h9678: y = 16'hfe00;
			16'h9679: y = 16'hfe00;
			16'h967a: y = 16'hfe00;
			16'h967b: y = 16'hfe00;
			16'h967c: y = 16'hfe00;
			16'h967d: y = 16'hfe00;
			16'h967e: y = 16'hfe00;
			16'h967f: y = 16'hfe00;
			16'h9680: y = 16'hfe00;
			16'h9681: y = 16'hfe00;
			16'h9682: y = 16'hfe00;
			16'h9683: y = 16'hfe00;
			16'h9684: y = 16'hfe00;
			16'h9685: y = 16'hfe00;
			16'h9686: y = 16'hfe00;
			16'h9687: y = 16'hfe00;
			16'h9688: y = 16'hfe00;
			16'h9689: y = 16'hfe00;
			16'h968a: y = 16'hfe00;
			16'h968b: y = 16'hfe00;
			16'h968c: y = 16'hfe00;
			16'h968d: y = 16'hfe00;
			16'h968e: y = 16'hfe00;
			16'h968f: y = 16'hfe00;
			16'h9690: y = 16'hfe00;
			16'h9691: y = 16'hfe00;
			16'h9692: y = 16'hfe00;
			16'h9693: y = 16'hfe00;
			16'h9694: y = 16'hfe00;
			16'h9695: y = 16'hfe00;
			16'h9696: y = 16'hfe00;
			16'h9697: y = 16'hfe00;
			16'h9698: y = 16'hfe00;
			16'h9699: y = 16'hfe00;
			16'h969a: y = 16'hfe00;
			16'h969b: y = 16'hfe00;
			16'h969c: y = 16'hfe00;
			16'h969d: y = 16'hfe00;
			16'h969e: y = 16'hfe00;
			16'h969f: y = 16'hfe00;
			16'h96a0: y = 16'hfe00;
			16'h96a1: y = 16'hfe00;
			16'h96a2: y = 16'hfe00;
			16'h96a3: y = 16'hfe00;
			16'h96a4: y = 16'hfe00;
			16'h96a5: y = 16'hfe00;
			16'h96a6: y = 16'hfe00;
			16'h96a7: y = 16'hfe00;
			16'h96a8: y = 16'hfe00;
			16'h96a9: y = 16'hfe00;
			16'h96aa: y = 16'hfe00;
			16'h96ab: y = 16'hfe00;
			16'h96ac: y = 16'hfe00;
			16'h96ad: y = 16'hfe00;
			16'h96ae: y = 16'hfe00;
			16'h96af: y = 16'hfe00;
			16'h96b0: y = 16'hfe00;
			16'h96b1: y = 16'hfe00;
			16'h96b2: y = 16'hfe00;
			16'h96b3: y = 16'hfe00;
			16'h96b4: y = 16'hfe00;
			16'h96b5: y = 16'hfe00;
			16'h96b6: y = 16'hfe00;
			16'h96b7: y = 16'hfe00;
			16'h96b8: y = 16'hfe00;
			16'h96b9: y = 16'hfe00;
			16'h96ba: y = 16'hfe00;
			16'h96bb: y = 16'hfe00;
			16'h96bc: y = 16'hfe00;
			16'h96bd: y = 16'hfe00;
			16'h96be: y = 16'hfe00;
			16'h96bf: y = 16'hfe00;
			16'h96c0: y = 16'hfe00;
			16'h96c1: y = 16'hfe00;
			16'h96c2: y = 16'hfe00;
			16'h96c3: y = 16'hfe00;
			16'h96c4: y = 16'hfe00;
			16'h96c5: y = 16'hfe00;
			16'h96c6: y = 16'hfe00;
			16'h96c7: y = 16'hfe00;
			16'h96c8: y = 16'hfe00;
			16'h96c9: y = 16'hfe00;
			16'h96ca: y = 16'hfe00;
			16'h96cb: y = 16'hfe00;
			16'h96cc: y = 16'hfe00;
			16'h96cd: y = 16'hfe00;
			16'h96ce: y = 16'hfe00;
			16'h96cf: y = 16'hfe00;
			16'h96d0: y = 16'hfe00;
			16'h96d1: y = 16'hfe00;
			16'h96d2: y = 16'hfe00;
			16'h96d3: y = 16'hfe00;
			16'h96d4: y = 16'hfe00;
			16'h96d5: y = 16'hfe00;
			16'h96d6: y = 16'hfe00;
			16'h96d7: y = 16'hfe00;
			16'h96d8: y = 16'hfe00;
			16'h96d9: y = 16'hfe00;
			16'h96da: y = 16'hfe00;
			16'h96db: y = 16'hfe00;
			16'h96dc: y = 16'hfe00;
			16'h96dd: y = 16'hfe00;
			16'h96de: y = 16'hfe00;
			16'h96df: y = 16'hfe00;
			16'h96e0: y = 16'hfe00;
			16'h96e1: y = 16'hfe00;
			16'h96e2: y = 16'hfe00;
			16'h96e3: y = 16'hfe00;
			16'h96e4: y = 16'hfe00;
			16'h96e5: y = 16'hfe00;
			16'h96e6: y = 16'hfe00;
			16'h96e7: y = 16'hfe00;
			16'h96e8: y = 16'hfe00;
			16'h96e9: y = 16'hfe00;
			16'h96ea: y = 16'hfe00;
			16'h96eb: y = 16'hfe00;
			16'h96ec: y = 16'hfe00;
			16'h96ed: y = 16'hfe00;
			16'h96ee: y = 16'hfe00;
			16'h96ef: y = 16'hfe00;
			16'h96f0: y = 16'hfe00;
			16'h96f1: y = 16'hfe00;
			16'h96f2: y = 16'hfe00;
			16'h96f3: y = 16'hfe00;
			16'h96f4: y = 16'hfe00;
			16'h96f5: y = 16'hfe00;
			16'h96f6: y = 16'hfe00;
			16'h96f7: y = 16'hfe00;
			16'h96f8: y = 16'hfe00;
			16'h96f9: y = 16'hfe00;
			16'h96fa: y = 16'hfe00;
			16'h96fb: y = 16'hfe00;
			16'h96fc: y = 16'hfe00;
			16'h96fd: y = 16'hfe00;
			16'h96fe: y = 16'hfe00;
			16'h96ff: y = 16'hfe00;
			16'h9700: y = 16'hfe00;
			16'h9701: y = 16'hfe00;
			16'h9702: y = 16'hfe00;
			16'h9703: y = 16'hfe00;
			16'h9704: y = 16'hfe00;
			16'h9705: y = 16'hfe00;
			16'h9706: y = 16'hfe00;
			16'h9707: y = 16'hfe00;
			16'h9708: y = 16'hfe00;
			16'h9709: y = 16'hfe00;
			16'h970a: y = 16'hfe00;
			16'h970b: y = 16'hfe00;
			16'h970c: y = 16'hfe00;
			16'h970d: y = 16'hfe00;
			16'h970e: y = 16'hfe00;
			16'h970f: y = 16'hfe00;
			16'h9710: y = 16'hfe00;
			16'h9711: y = 16'hfe00;
			16'h9712: y = 16'hfe00;
			16'h9713: y = 16'hfe00;
			16'h9714: y = 16'hfe00;
			16'h9715: y = 16'hfe00;
			16'h9716: y = 16'hfe00;
			16'h9717: y = 16'hfe00;
			16'h9718: y = 16'hfe00;
			16'h9719: y = 16'hfe00;
			16'h971a: y = 16'hfe00;
			16'h971b: y = 16'hfe00;
			16'h971c: y = 16'hfe00;
			16'h971d: y = 16'hfe00;
			16'h971e: y = 16'hfe00;
			16'h971f: y = 16'hfe00;
			16'h9720: y = 16'hfe00;
			16'h9721: y = 16'hfe00;
			16'h9722: y = 16'hfe00;
			16'h9723: y = 16'hfe00;
			16'h9724: y = 16'hfe00;
			16'h9725: y = 16'hfe00;
			16'h9726: y = 16'hfe00;
			16'h9727: y = 16'hfe00;
			16'h9728: y = 16'hfe00;
			16'h9729: y = 16'hfe00;
			16'h972a: y = 16'hfe00;
			16'h972b: y = 16'hfe00;
			16'h972c: y = 16'hfe00;
			16'h972d: y = 16'hfe00;
			16'h972e: y = 16'hfe00;
			16'h972f: y = 16'hfe00;
			16'h9730: y = 16'hfe00;
			16'h9731: y = 16'hfe00;
			16'h9732: y = 16'hfe00;
			16'h9733: y = 16'hfe00;
			16'h9734: y = 16'hfe00;
			16'h9735: y = 16'hfe00;
			16'h9736: y = 16'hfe00;
			16'h9737: y = 16'hfe00;
			16'h9738: y = 16'hfe00;
			16'h9739: y = 16'hfe00;
			16'h973a: y = 16'hfe00;
			16'h973b: y = 16'hfe00;
			16'h973c: y = 16'hfe00;
			16'h973d: y = 16'hfe00;
			16'h973e: y = 16'hfe00;
			16'h973f: y = 16'hfe00;
			16'h9740: y = 16'hfe00;
			16'h9741: y = 16'hfe00;
			16'h9742: y = 16'hfe00;
			16'h9743: y = 16'hfe00;
			16'h9744: y = 16'hfe00;
			16'h9745: y = 16'hfe00;
			16'h9746: y = 16'hfe00;
			16'h9747: y = 16'hfe00;
			16'h9748: y = 16'hfe00;
			16'h9749: y = 16'hfe00;
			16'h974a: y = 16'hfe00;
			16'h974b: y = 16'hfe00;
			16'h974c: y = 16'hfe00;
			16'h974d: y = 16'hfe00;
			16'h974e: y = 16'hfe00;
			16'h974f: y = 16'hfe00;
			16'h9750: y = 16'hfe00;
			16'h9751: y = 16'hfe00;
			16'h9752: y = 16'hfe00;
			16'h9753: y = 16'hfe00;
			16'h9754: y = 16'hfe00;
			16'h9755: y = 16'hfe00;
			16'h9756: y = 16'hfe00;
			16'h9757: y = 16'hfe00;
			16'h9758: y = 16'hfe00;
			16'h9759: y = 16'hfe00;
			16'h975a: y = 16'hfe00;
			16'h975b: y = 16'hfe00;
			16'h975c: y = 16'hfe00;
			16'h975d: y = 16'hfe00;
			16'h975e: y = 16'hfe00;
			16'h975f: y = 16'hfe00;
			16'h9760: y = 16'hfe00;
			16'h9761: y = 16'hfe00;
			16'h9762: y = 16'hfe00;
			16'h9763: y = 16'hfe00;
			16'h9764: y = 16'hfe00;
			16'h9765: y = 16'hfe00;
			16'h9766: y = 16'hfe00;
			16'h9767: y = 16'hfe00;
			16'h9768: y = 16'hfe00;
			16'h9769: y = 16'hfe00;
			16'h976a: y = 16'hfe00;
			16'h976b: y = 16'hfe00;
			16'h976c: y = 16'hfe00;
			16'h976d: y = 16'hfe00;
			16'h976e: y = 16'hfe00;
			16'h976f: y = 16'hfe00;
			16'h9770: y = 16'hfe00;
			16'h9771: y = 16'hfe00;
			16'h9772: y = 16'hfe00;
			16'h9773: y = 16'hfe00;
			16'h9774: y = 16'hfe00;
			16'h9775: y = 16'hfe00;
			16'h9776: y = 16'hfe00;
			16'h9777: y = 16'hfe00;
			16'h9778: y = 16'hfe00;
			16'h9779: y = 16'hfe00;
			16'h977a: y = 16'hfe00;
			16'h977b: y = 16'hfe00;
			16'h977c: y = 16'hfe00;
			16'h977d: y = 16'hfe00;
			16'h977e: y = 16'hfe00;
			16'h977f: y = 16'hfe00;
			16'h9780: y = 16'hfe00;
			16'h9781: y = 16'hfe00;
			16'h9782: y = 16'hfe00;
			16'h9783: y = 16'hfe00;
			16'h9784: y = 16'hfe00;
			16'h9785: y = 16'hfe00;
			16'h9786: y = 16'hfe00;
			16'h9787: y = 16'hfe00;
			16'h9788: y = 16'hfe00;
			16'h9789: y = 16'hfe00;
			16'h978a: y = 16'hfe00;
			16'h978b: y = 16'hfe00;
			16'h978c: y = 16'hfe00;
			16'h978d: y = 16'hfe00;
			16'h978e: y = 16'hfe00;
			16'h978f: y = 16'hfe00;
			16'h9790: y = 16'hfe00;
			16'h9791: y = 16'hfe00;
			16'h9792: y = 16'hfe00;
			16'h9793: y = 16'hfe00;
			16'h9794: y = 16'hfe00;
			16'h9795: y = 16'hfe00;
			16'h9796: y = 16'hfe00;
			16'h9797: y = 16'hfe00;
			16'h9798: y = 16'hfe00;
			16'h9799: y = 16'hfe00;
			16'h979a: y = 16'hfe00;
			16'h979b: y = 16'hfe00;
			16'h979c: y = 16'hfe00;
			16'h979d: y = 16'hfe00;
			16'h979e: y = 16'hfe00;
			16'h979f: y = 16'hfe00;
			16'h97a0: y = 16'hfe00;
			16'h97a1: y = 16'hfe00;
			16'h97a2: y = 16'hfe00;
			16'h97a3: y = 16'hfe00;
			16'h97a4: y = 16'hfe00;
			16'h97a5: y = 16'hfe00;
			16'h97a6: y = 16'hfe00;
			16'h97a7: y = 16'hfe00;
			16'h97a8: y = 16'hfe00;
			16'h97a9: y = 16'hfe00;
			16'h97aa: y = 16'hfe00;
			16'h97ab: y = 16'hfe00;
			16'h97ac: y = 16'hfe00;
			16'h97ad: y = 16'hfe00;
			16'h97ae: y = 16'hfe00;
			16'h97af: y = 16'hfe00;
			16'h97b0: y = 16'hfe00;
			16'h97b1: y = 16'hfe00;
			16'h97b2: y = 16'hfe00;
			16'h97b3: y = 16'hfe00;
			16'h97b4: y = 16'hfe00;
			16'h97b5: y = 16'hfe00;
			16'h97b6: y = 16'hfe00;
			16'h97b7: y = 16'hfe00;
			16'h97b8: y = 16'hfe00;
			16'h97b9: y = 16'hfe00;
			16'h97ba: y = 16'hfe00;
			16'h97bb: y = 16'hfe00;
			16'h97bc: y = 16'hfe00;
			16'h97bd: y = 16'hfe00;
			16'h97be: y = 16'hfe00;
			16'h97bf: y = 16'hfe00;
			16'h97c0: y = 16'hfe00;
			16'h97c1: y = 16'hfe00;
			16'h97c2: y = 16'hfe00;
			16'h97c3: y = 16'hfe00;
			16'h97c4: y = 16'hfe00;
			16'h97c5: y = 16'hfe00;
			16'h97c6: y = 16'hfe00;
			16'h97c7: y = 16'hfe00;
			16'h97c8: y = 16'hfe00;
			16'h97c9: y = 16'hfe00;
			16'h97ca: y = 16'hfe00;
			16'h97cb: y = 16'hfe00;
			16'h97cc: y = 16'hfe00;
			16'h97cd: y = 16'hfe00;
			16'h97ce: y = 16'hfe00;
			16'h97cf: y = 16'hfe00;
			16'h97d0: y = 16'hfe00;
			16'h97d1: y = 16'hfe00;
			16'h97d2: y = 16'hfe00;
			16'h97d3: y = 16'hfe00;
			16'h97d4: y = 16'hfe00;
			16'h97d5: y = 16'hfe00;
			16'h97d6: y = 16'hfe00;
			16'h97d7: y = 16'hfe00;
			16'h97d8: y = 16'hfe00;
			16'h97d9: y = 16'hfe00;
			16'h97da: y = 16'hfe00;
			16'h97db: y = 16'hfe00;
			16'h97dc: y = 16'hfe00;
			16'h97dd: y = 16'hfe00;
			16'h97de: y = 16'hfe00;
			16'h97df: y = 16'hfe00;
			16'h97e0: y = 16'hfe00;
			16'h97e1: y = 16'hfe00;
			16'h97e2: y = 16'hfe00;
			16'h97e3: y = 16'hfe00;
			16'h97e4: y = 16'hfe00;
			16'h97e5: y = 16'hfe00;
			16'h97e6: y = 16'hfe00;
			16'h97e7: y = 16'hfe00;
			16'h97e8: y = 16'hfe00;
			16'h97e9: y = 16'hfe00;
			16'h97ea: y = 16'hfe00;
			16'h97eb: y = 16'hfe00;
			16'h97ec: y = 16'hfe00;
			16'h97ed: y = 16'hfe00;
			16'h97ee: y = 16'hfe00;
			16'h97ef: y = 16'hfe00;
			16'h97f0: y = 16'hfe00;
			16'h97f1: y = 16'hfe00;
			16'h97f2: y = 16'hfe00;
			16'h97f3: y = 16'hfe00;
			16'h97f4: y = 16'hfe00;
			16'h97f5: y = 16'hfe00;
			16'h97f6: y = 16'hfe00;
			16'h97f7: y = 16'hfe00;
			16'h97f8: y = 16'hfe00;
			16'h97f9: y = 16'hfe00;
			16'h97fa: y = 16'hfe00;
			16'h97fb: y = 16'hfe00;
			16'h97fc: y = 16'hfe00;
			16'h97fd: y = 16'hfe00;
			16'h97fe: y = 16'hfe00;
			16'h97ff: y = 16'hfe00;
			16'h9800: y = 16'hfe00;
			16'h9801: y = 16'hfe00;
			16'h9802: y = 16'hfe00;
			16'h9803: y = 16'hfe00;
			16'h9804: y = 16'hfe00;
			16'h9805: y = 16'hfe00;
			16'h9806: y = 16'hfe00;
			16'h9807: y = 16'hfe00;
			16'h9808: y = 16'hfe00;
			16'h9809: y = 16'hfe00;
			16'h980a: y = 16'hfe00;
			16'h980b: y = 16'hfe00;
			16'h980c: y = 16'hfe00;
			16'h980d: y = 16'hfe00;
			16'h980e: y = 16'hfe00;
			16'h980f: y = 16'hfe00;
			16'h9810: y = 16'hfe00;
			16'h9811: y = 16'hfe00;
			16'h9812: y = 16'hfe00;
			16'h9813: y = 16'hfe00;
			16'h9814: y = 16'hfe00;
			16'h9815: y = 16'hfe00;
			16'h9816: y = 16'hfe00;
			16'h9817: y = 16'hfe00;
			16'h9818: y = 16'hfe00;
			16'h9819: y = 16'hfe00;
			16'h981a: y = 16'hfe00;
			16'h981b: y = 16'hfe00;
			16'h981c: y = 16'hfe00;
			16'h981d: y = 16'hfe00;
			16'h981e: y = 16'hfe00;
			16'h981f: y = 16'hfe00;
			16'h9820: y = 16'hfe00;
			16'h9821: y = 16'hfe00;
			16'h9822: y = 16'hfe00;
			16'h9823: y = 16'hfe00;
			16'h9824: y = 16'hfe00;
			16'h9825: y = 16'hfe00;
			16'h9826: y = 16'hfe00;
			16'h9827: y = 16'hfe00;
			16'h9828: y = 16'hfe00;
			16'h9829: y = 16'hfe00;
			16'h982a: y = 16'hfe00;
			16'h982b: y = 16'hfe00;
			16'h982c: y = 16'hfe00;
			16'h982d: y = 16'hfe00;
			16'h982e: y = 16'hfe00;
			16'h982f: y = 16'hfe00;
			16'h9830: y = 16'hfe00;
			16'h9831: y = 16'hfe00;
			16'h9832: y = 16'hfe00;
			16'h9833: y = 16'hfe00;
			16'h9834: y = 16'hfe00;
			16'h9835: y = 16'hfe00;
			16'h9836: y = 16'hfe00;
			16'h9837: y = 16'hfe00;
			16'h9838: y = 16'hfe00;
			16'h9839: y = 16'hfe00;
			16'h983a: y = 16'hfe00;
			16'h983b: y = 16'hfe00;
			16'h983c: y = 16'hfe00;
			16'h983d: y = 16'hfe00;
			16'h983e: y = 16'hfe00;
			16'h983f: y = 16'hfe00;
			16'h9840: y = 16'hfe00;
			16'h9841: y = 16'hfe00;
			16'h9842: y = 16'hfe00;
			16'h9843: y = 16'hfe00;
			16'h9844: y = 16'hfe00;
			16'h9845: y = 16'hfe00;
			16'h9846: y = 16'hfe00;
			16'h9847: y = 16'hfe00;
			16'h9848: y = 16'hfe00;
			16'h9849: y = 16'hfe00;
			16'h984a: y = 16'hfe00;
			16'h984b: y = 16'hfe00;
			16'h984c: y = 16'hfe00;
			16'h984d: y = 16'hfe00;
			16'h984e: y = 16'hfe00;
			16'h984f: y = 16'hfe00;
			16'h9850: y = 16'hfe00;
			16'h9851: y = 16'hfe00;
			16'h9852: y = 16'hfe00;
			16'h9853: y = 16'hfe00;
			16'h9854: y = 16'hfe00;
			16'h9855: y = 16'hfe00;
			16'h9856: y = 16'hfe00;
			16'h9857: y = 16'hfe00;
			16'h9858: y = 16'hfe00;
			16'h9859: y = 16'hfe00;
			16'h985a: y = 16'hfe00;
			16'h985b: y = 16'hfe00;
			16'h985c: y = 16'hfe00;
			16'h985d: y = 16'hfe00;
			16'h985e: y = 16'hfe00;
			16'h985f: y = 16'hfe00;
			16'h9860: y = 16'hfe00;
			16'h9861: y = 16'hfe00;
			16'h9862: y = 16'hfe00;
			16'h9863: y = 16'hfe00;
			16'h9864: y = 16'hfe00;
			16'h9865: y = 16'hfe00;
			16'h9866: y = 16'hfe00;
			16'h9867: y = 16'hfe00;
			16'h9868: y = 16'hfe00;
			16'h9869: y = 16'hfe00;
			16'h986a: y = 16'hfe00;
			16'h986b: y = 16'hfe00;
			16'h986c: y = 16'hfe00;
			16'h986d: y = 16'hfe00;
			16'h986e: y = 16'hfe00;
			16'h986f: y = 16'hfe00;
			16'h9870: y = 16'hfe00;
			16'h9871: y = 16'hfe00;
			16'h9872: y = 16'hfe00;
			16'h9873: y = 16'hfe00;
			16'h9874: y = 16'hfe00;
			16'h9875: y = 16'hfe00;
			16'h9876: y = 16'hfe00;
			16'h9877: y = 16'hfe00;
			16'h9878: y = 16'hfe00;
			16'h9879: y = 16'hfe00;
			16'h987a: y = 16'hfe00;
			16'h987b: y = 16'hfe00;
			16'h987c: y = 16'hfe00;
			16'h987d: y = 16'hfe00;
			16'h987e: y = 16'hfe00;
			16'h987f: y = 16'hfe00;
			16'h9880: y = 16'hfe00;
			16'h9881: y = 16'hfe00;
			16'h9882: y = 16'hfe00;
			16'h9883: y = 16'hfe00;
			16'h9884: y = 16'hfe00;
			16'h9885: y = 16'hfe00;
			16'h9886: y = 16'hfe00;
			16'h9887: y = 16'hfe00;
			16'h9888: y = 16'hfe00;
			16'h9889: y = 16'hfe00;
			16'h988a: y = 16'hfe00;
			16'h988b: y = 16'hfe00;
			16'h988c: y = 16'hfe00;
			16'h988d: y = 16'hfe00;
			16'h988e: y = 16'hfe00;
			16'h988f: y = 16'hfe00;
			16'h9890: y = 16'hfe00;
			16'h9891: y = 16'hfe00;
			16'h9892: y = 16'hfe00;
			16'h9893: y = 16'hfe00;
			16'h9894: y = 16'hfe00;
			16'h9895: y = 16'hfe00;
			16'h9896: y = 16'hfe00;
			16'h9897: y = 16'hfe00;
			16'h9898: y = 16'hfe00;
			16'h9899: y = 16'hfe00;
			16'h989a: y = 16'hfe00;
			16'h989b: y = 16'hfe00;
			16'h989c: y = 16'hfe00;
			16'h989d: y = 16'hfe00;
			16'h989e: y = 16'hfe00;
			16'h989f: y = 16'hfe00;
			16'h98a0: y = 16'hfe00;
			16'h98a1: y = 16'hfe00;
			16'h98a2: y = 16'hfe00;
			16'h98a3: y = 16'hfe00;
			16'h98a4: y = 16'hfe00;
			16'h98a5: y = 16'hfe00;
			16'h98a6: y = 16'hfe00;
			16'h98a7: y = 16'hfe00;
			16'h98a8: y = 16'hfe00;
			16'h98a9: y = 16'hfe00;
			16'h98aa: y = 16'hfe00;
			16'h98ab: y = 16'hfe00;
			16'h98ac: y = 16'hfe00;
			16'h98ad: y = 16'hfe00;
			16'h98ae: y = 16'hfe00;
			16'h98af: y = 16'hfe00;
			16'h98b0: y = 16'hfe00;
			16'h98b1: y = 16'hfe00;
			16'h98b2: y = 16'hfe00;
			16'h98b3: y = 16'hfe00;
			16'h98b4: y = 16'hfe00;
			16'h98b5: y = 16'hfe00;
			16'h98b6: y = 16'hfe00;
			16'h98b7: y = 16'hfe00;
			16'h98b8: y = 16'hfe00;
			16'h98b9: y = 16'hfe00;
			16'h98ba: y = 16'hfe00;
			16'h98bb: y = 16'hfe00;
			16'h98bc: y = 16'hfe00;
			16'h98bd: y = 16'hfe00;
			16'h98be: y = 16'hfe00;
			16'h98bf: y = 16'hfe00;
			16'h98c0: y = 16'hfe00;
			16'h98c1: y = 16'hfe00;
			16'h98c2: y = 16'hfe00;
			16'h98c3: y = 16'hfe00;
			16'h98c4: y = 16'hfe00;
			16'h98c5: y = 16'hfe00;
			16'h98c6: y = 16'hfe00;
			16'h98c7: y = 16'hfe00;
			16'h98c8: y = 16'hfe00;
			16'h98c9: y = 16'hfe00;
			16'h98ca: y = 16'hfe00;
			16'h98cb: y = 16'hfe00;
			16'h98cc: y = 16'hfe00;
			16'h98cd: y = 16'hfe00;
			16'h98ce: y = 16'hfe00;
			16'h98cf: y = 16'hfe00;
			16'h98d0: y = 16'hfe00;
			16'h98d1: y = 16'hfe00;
			16'h98d2: y = 16'hfe00;
			16'h98d3: y = 16'hfe00;
			16'h98d4: y = 16'hfe00;
			16'h98d5: y = 16'hfe00;
			16'h98d6: y = 16'hfe00;
			16'h98d7: y = 16'hfe00;
			16'h98d8: y = 16'hfe00;
			16'h98d9: y = 16'hfe00;
			16'h98da: y = 16'hfe00;
			16'h98db: y = 16'hfe00;
			16'h98dc: y = 16'hfe00;
			16'h98dd: y = 16'hfe00;
			16'h98de: y = 16'hfe00;
			16'h98df: y = 16'hfe00;
			16'h98e0: y = 16'hfe00;
			16'h98e1: y = 16'hfe00;
			16'h98e2: y = 16'hfe00;
			16'h98e3: y = 16'hfe00;
			16'h98e4: y = 16'hfe00;
			16'h98e5: y = 16'hfe00;
			16'h98e6: y = 16'hfe00;
			16'h98e7: y = 16'hfe00;
			16'h98e8: y = 16'hfe00;
			16'h98e9: y = 16'hfe00;
			16'h98ea: y = 16'hfe00;
			16'h98eb: y = 16'hfe00;
			16'h98ec: y = 16'hfe00;
			16'h98ed: y = 16'hfe00;
			16'h98ee: y = 16'hfe00;
			16'h98ef: y = 16'hfe00;
			16'h98f0: y = 16'hfe00;
			16'h98f1: y = 16'hfe00;
			16'h98f2: y = 16'hfe00;
			16'h98f3: y = 16'hfe00;
			16'h98f4: y = 16'hfe00;
			16'h98f5: y = 16'hfe00;
			16'h98f6: y = 16'hfe00;
			16'h98f7: y = 16'hfe00;
			16'h98f8: y = 16'hfe00;
			16'h98f9: y = 16'hfe00;
			16'h98fa: y = 16'hfe00;
			16'h98fb: y = 16'hfe00;
			16'h98fc: y = 16'hfe00;
			16'h98fd: y = 16'hfe00;
			16'h98fe: y = 16'hfe00;
			16'h98ff: y = 16'hfe00;
			16'h9900: y = 16'hfe00;
			16'h9901: y = 16'hfe00;
			16'h9902: y = 16'hfe00;
			16'h9903: y = 16'hfe00;
			16'h9904: y = 16'hfe00;
			16'h9905: y = 16'hfe00;
			16'h9906: y = 16'hfe00;
			16'h9907: y = 16'hfe00;
			16'h9908: y = 16'hfe00;
			16'h9909: y = 16'hfe00;
			16'h990a: y = 16'hfe00;
			16'h990b: y = 16'hfe00;
			16'h990c: y = 16'hfe00;
			16'h990d: y = 16'hfe00;
			16'h990e: y = 16'hfe00;
			16'h990f: y = 16'hfe00;
			16'h9910: y = 16'hfe00;
			16'h9911: y = 16'hfe00;
			16'h9912: y = 16'hfe00;
			16'h9913: y = 16'hfe00;
			16'h9914: y = 16'hfe00;
			16'h9915: y = 16'hfe00;
			16'h9916: y = 16'hfe00;
			16'h9917: y = 16'hfe00;
			16'h9918: y = 16'hfe00;
			16'h9919: y = 16'hfe00;
			16'h991a: y = 16'hfe00;
			16'h991b: y = 16'hfe00;
			16'h991c: y = 16'hfe00;
			16'h991d: y = 16'hfe00;
			16'h991e: y = 16'hfe00;
			16'h991f: y = 16'hfe00;
			16'h9920: y = 16'hfe00;
			16'h9921: y = 16'hfe00;
			16'h9922: y = 16'hfe00;
			16'h9923: y = 16'hfe00;
			16'h9924: y = 16'hfe00;
			16'h9925: y = 16'hfe00;
			16'h9926: y = 16'hfe00;
			16'h9927: y = 16'hfe00;
			16'h9928: y = 16'hfe00;
			16'h9929: y = 16'hfe00;
			16'h992a: y = 16'hfe00;
			16'h992b: y = 16'hfe00;
			16'h992c: y = 16'hfe00;
			16'h992d: y = 16'hfe00;
			16'h992e: y = 16'hfe00;
			16'h992f: y = 16'hfe00;
			16'h9930: y = 16'hfe00;
			16'h9931: y = 16'hfe00;
			16'h9932: y = 16'hfe00;
			16'h9933: y = 16'hfe00;
			16'h9934: y = 16'hfe00;
			16'h9935: y = 16'hfe00;
			16'h9936: y = 16'hfe00;
			16'h9937: y = 16'hfe00;
			16'h9938: y = 16'hfe00;
			16'h9939: y = 16'hfe00;
			16'h993a: y = 16'hfe00;
			16'h993b: y = 16'hfe00;
			16'h993c: y = 16'hfe00;
			16'h993d: y = 16'hfe00;
			16'h993e: y = 16'hfe00;
			16'h993f: y = 16'hfe00;
			16'h9940: y = 16'hfe00;
			16'h9941: y = 16'hfe00;
			16'h9942: y = 16'hfe00;
			16'h9943: y = 16'hfe00;
			16'h9944: y = 16'hfe00;
			16'h9945: y = 16'hfe00;
			16'h9946: y = 16'hfe00;
			16'h9947: y = 16'hfe00;
			16'h9948: y = 16'hfe00;
			16'h9949: y = 16'hfe00;
			16'h994a: y = 16'hfe00;
			16'h994b: y = 16'hfe00;
			16'h994c: y = 16'hfe00;
			16'h994d: y = 16'hfe00;
			16'h994e: y = 16'hfe00;
			16'h994f: y = 16'hfe00;
			16'h9950: y = 16'hfe00;
			16'h9951: y = 16'hfe00;
			16'h9952: y = 16'hfe00;
			16'h9953: y = 16'hfe00;
			16'h9954: y = 16'hfe00;
			16'h9955: y = 16'hfe00;
			16'h9956: y = 16'hfe00;
			16'h9957: y = 16'hfe00;
			16'h9958: y = 16'hfe00;
			16'h9959: y = 16'hfe00;
			16'h995a: y = 16'hfe00;
			16'h995b: y = 16'hfe00;
			16'h995c: y = 16'hfe00;
			16'h995d: y = 16'hfe00;
			16'h995e: y = 16'hfe00;
			16'h995f: y = 16'hfe00;
			16'h9960: y = 16'hfe00;
			16'h9961: y = 16'hfe00;
			16'h9962: y = 16'hfe00;
			16'h9963: y = 16'hfe00;
			16'h9964: y = 16'hfe00;
			16'h9965: y = 16'hfe00;
			16'h9966: y = 16'hfe00;
			16'h9967: y = 16'hfe00;
			16'h9968: y = 16'hfe00;
			16'h9969: y = 16'hfe00;
			16'h996a: y = 16'hfe00;
			16'h996b: y = 16'hfe00;
			16'h996c: y = 16'hfe00;
			16'h996d: y = 16'hfe00;
			16'h996e: y = 16'hfe00;
			16'h996f: y = 16'hfe00;
			16'h9970: y = 16'hfe00;
			16'h9971: y = 16'hfe00;
			16'h9972: y = 16'hfe00;
			16'h9973: y = 16'hfe00;
			16'h9974: y = 16'hfe00;
			16'h9975: y = 16'hfe00;
			16'h9976: y = 16'hfe00;
			16'h9977: y = 16'hfe00;
			16'h9978: y = 16'hfe00;
			16'h9979: y = 16'hfe00;
			16'h997a: y = 16'hfe00;
			16'h997b: y = 16'hfe00;
			16'h997c: y = 16'hfe00;
			16'h997d: y = 16'hfe00;
			16'h997e: y = 16'hfe00;
			16'h997f: y = 16'hfe00;
			16'h9980: y = 16'hfe00;
			16'h9981: y = 16'hfe00;
			16'h9982: y = 16'hfe00;
			16'h9983: y = 16'hfe00;
			16'h9984: y = 16'hfe00;
			16'h9985: y = 16'hfe00;
			16'h9986: y = 16'hfe00;
			16'h9987: y = 16'hfe00;
			16'h9988: y = 16'hfe00;
			16'h9989: y = 16'hfe00;
			16'h998a: y = 16'hfe00;
			16'h998b: y = 16'hfe00;
			16'h998c: y = 16'hfe00;
			16'h998d: y = 16'hfe00;
			16'h998e: y = 16'hfe00;
			16'h998f: y = 16'hfe00;
			16'h9990: y = 16'hfe00;
			16'h9991: y = 16'hfe00;
			16'h9992: y = 16'hfe00;
			16'h9993: y = 16'hfe00;
			16'h9994: y = 16'hfe00;
			16'h9995: y = 16'hfe00;
			16'h9996: y = 16'hfe00;
			16'h9997: y = 16'hfe00;
			16'h9998: y = 16'hfe00;
			16'h9999: y = 16'hfe00;
			16'h999a: y = 16'hfe00;
			16'h999b: y = 16'hfe00;
			16'h999c: y = 16'hfe00;
			16'h999d: y = 16'hfe00;
			16'h999e: y = 16'hfe00;
			16'h999f: y = 16'hfe00;
			16'h99a0: y = 16'hfe00;
			16'h99a1: y = 16'hfe00;
			16'h99a2: y = 16'hfe00;
			16'h99a3: y = 16'hfe00;
			16'h99a4: y = 16'hfe00;
			16'h99a5: y = 16'hfe00;
			16'h99a6: y = 16'hfe00;
			16'h99a7: y = 16'hfe00;
			16'h99a8: y = 16'hfe00;
			16'h99a9: y = 16'hfe00;
			16'h99aa: y = 16'hfe00;
			16'h99ab: y = 16'hfe00;
			16'h99ac: y = 16'hfe00;
			16'h99ad: y = 16'hfe00;
			16'h99ae: y = 16'hfe00;
			16'h99af: y = 16'hfe00;
			16'h99b0: y = 16'hfe00;
			16'h99b1: y = 16'hfe00;
			16'h99b2: y = 16'hfe00;
			16'h99b3: y = 16'hfe00;
			16'h99b4: y = 16'hfe00;
			16'h99b5: y = 16'hfe00;
			16'h99b6: y = 16'hfe00;
			16'h99b7: y = 16'hfe00;
			16'h99b8: y = 16'hfe00;
			16'h99b9: y = 16'hfe00;
			16'h99ba: y = 16'hfe00;
			16'h99bb: y = 16'hfe00;
			16'h99bc: y = 16'hfe00;
			16'h99bd: y = 16'hfe00;
			16'h99be: y = 16'hfe00;
			16'h99bf: y = 16'hfe00;
			16'h99c0: y = 16'hfe00;
			16'h99c1: y = 16'hfe00;
			16'h99c2: y = 16'hfe00;
			16'h99c3: y = 16'hfe00;
			16'h99c4: y = 16'hfe00;
			16'h99c5: y = 16'hfe00;
			16'h99c6: y = 16'hfe00;
			16'h99c7: y = 16'hfe00;
			16'h99c8: y = 16'hfe00;
			16'h99c9: y = 16'hfe00;
			16'h99ca: y = 16'hfe00;
			16'h99cb: y = 16'hfe00;
			16'h99cc: y = 16'hfe00;
			16'h99cd: y = 16'hfe00;
			16'h99ce: y = 16'hfe00;
			16'h99cf: y = 16'hfe00;
			16'h99d0: y = 16'hfe00;
			16'h99d1: y = 16'hfe00;
			16'h99d2: y = 16'hfe00;
			16'h99d3: y = 16'hfe00;
			16'h99d4: y = 16'hfe00;
			16'h99d5: y = 16'hfe00;
			16'h99d6: y = 16'hfe00;
			16'h99d7: y = 16'hfe00;
			16'h99d8: y = 16'hfe00;
			16'h99d9: y = 16'hfe00;
			16'h99da: y = 16'hfe00;
			16'h99db: y = 16'hfe00;
			16'h99dc: y = 16'hfe00;
			16'h99dd: y = 16'hfe00;
			16'h99de: y = 16'hfe00;
			16'h99df: y = 16'hfe00;
			16'h99e0: y = 16'hfe00;
			16'h99e1: y = 16'hfe00;
			16'h99e2: y = 16'hfe00;
			16'h99e3: y = 16'hfe00;
			16'h99e4: y = 16'hfe00;
			16'h99e5: y = 16'hfe00;
			16'h99e6: y = 16'hfe00;
			16'h99e7: y = 16'hfe00;
			16'h99e8: y = 16'hfe00;
			16'h99e9: y = 16'hfe00;
			16'h99ea: y = 16'hfe00;
			16'h99eb: y = 16'hfe00;
			16'h99ec: y = 16'hfe00;
			16'h99ed: y = 16'hfe00;
			16'h99ee: y = 16'hfe00;
			16'h99ef: y = 16'hfe00;
			16'h99f0: y = 16'hfe00;
			16'h99f1: y = 16'hfe00;
			16'h99f2: y = 16'hfe00;
			16'h99f3: y = 16'hfe00;
			16'h99f4: y = 16'hfe00;
			16'h99f5: y = 16'hfe00;
			16'h99f6: y = 16'hfe00;
			16'h99f7: y = 16'hfe00;
			16'h99f8: y = 16'hfe00;
			16'h99f9: y = 16'hfe00;
			16'h99fa: y = 16'hfe00;
			16'h99fb: y = 16'hfe00;
			16'h99fc: y = 16'hfe00;
			16'h99fd: y = 16'hfe00;
			16'h99fe: y = 16'hfe00;
			16'h99ff: y = 16'hfe00;
			16'h9a00: y = 16'hfe00;
			16'h9a01: y = 16'hfe00;
			16'h9a02: y = 16'hfe00;
			16'h9a03: y = 16'hfe00;
			16'h9a04: y = 16'hfe00;
			16'h9a05: y = 16'hfe00;
			16'h9a06: y = 16'hfe00;
			16'h9a07: y = 16'hfe00;
			16'h9a08: y = 16'hfe00;
			16'h9a09: y = 16'hfe00;
			16'h9a0a: y = 16'hfe00;
			16'h9a0b: y = 16'hfe00;
			16'h9a0c: y = 16'hfe00;
			16'h9a0d: y = 16'hfe00;
			16'h9a0e: y = 16'hfe00;
			16'h9a0f: y = 16'hfe00;
			16'h9a10: y = 16'hfe00;
			16'h9a11: y = 16'hfe00;
			16'h9a12: y = 16'hfe00;
			16'h9a13: y = 16'hfe00;
			16'h9a14: y = 16'hfe00;
			16'h9a15: y = 16'hfe00;
			16'h9a16: y = 16'hfe00;
			16'h9a17: y = 16'hfe00;
			16'h9a18: y = 16'hfe00;
			16'h9a19: y = 16'hfe00;
			16'h9a1a: y = 16'hfe00;
			16'h9a1b: y = 16'hfe00;
			16'h9a1c: y = 16'hfe00;
			16'h9a1d: y = 16'hfe00;
			16'h9a1e: y = 16'hfe00;
			16'h9a1f: y = 16'hfe00;
			16'h9a20: y = 16'hfe00;
			16'h9a21: y = 16'hfe00;
			16'h9a22: y = 16'hfe00;
			16'h9a23: y = 16'hfe00;
			16'h9a24: y = 16'hfe00;
			16'h9a25: y = 16'hfe00;
			16'h9a26: y = 16'hfe00;
			16'h9a27: y = 16'hfe00;
			16'h9a28: y = 16'hfe00;
			16'h9a29: y = 16'hfe00;
			16'h9a2a: y = 16'hfe00;
			16'h9a2b: y = 16'hfe00;
			16'h9a2c: y = 16'hfe00;
			16'h9a2d: y = 16'hfe00;
			16'h9a2e: y = 16'hfe00;
			16'h9a2f: y = 16'hfe00;
			16'h9a30: y = 16'hfe00;
			16'h9a31: y = 16'hfe00;
			16'h9a32: y = 16'hfe00;
			16'h9a33: y = 16'hfe00;
			16'h9a34: y = 16'hfe00;
			16'h9a35: y = 16'hfe00;
			16'h9a36: y = 16'hfe00;
			16'h9a37: y = 16'hfe00;
			16'h9a38: y = 16'hfe00;
			16'h9a39: y = 16'hfe00;
			16'h9a3a: y = 16'hfe00;
			16'h9a3b: y = 16'hfe00;
			16'h9a3c: y = 16'hfe00;
			16'h9a3d: y = 16'hfe00;
			16'h9a3e: y = 16'hfe00;
			16'h9a3f: y = 16'hfe00;
			16'h9a40: y = 16'hfe00;
			16'h9a41: y = 16'hfe00;
			16'h9a42: y = 16'hfe00;
			16'h9a43: y = 16'hfe00;
			16'h9a44: y = 16'hfe00;
			16'h9a45: y = 16'hfe00;
			16'h9a46: y = 16'hfe00;
			16'h9a47: y = 16'hfe00;
			16'h9a48: y = 16'hfe00;
			16'h9a49: y = 16'hfe00;
			16'h9a4a: y = 16'hfe00;
			16'h9a4b: y = 16'hfe00;
			16'h9a4c: y = 16'hfe00;
			16'h9a4d: y = 16'hfe00;
			16'h9a4e: y = 16'hfe00;
			16'h9a4f: y = 16'hfe00;
			16'h9a50: y = 16'hfe00;
			16'h9a51: y = 16'hfe00;
			16'h9a52: y = 16'hfe00;
			16'h9a53: y = 16'hfe00;
			16'h9a54: y = 16'hfe00;
			16'h9a55: y = 16'hfe00;
			16'h9a56: y = 16'hfe00;
			16'h9a57: y = 16'hfe00;
			16'h9a58: y = 16'hfe00;
			16'h9a59: y = 16'hfe00;
			16'h9a5a: y = 16'hfe00;
			16'h9a5b: y = 16'hfe00;
			16'h9a5c: y = 16'hfe00;
			16'h9a5d: y = 16'hfe00;
			16'h9a5e: y = 16'hfe00;
			16'h9a5f: y = 16'hfe00;
			16'h9a60: y = 16'hfe00;
			16'h9a61: y = 16'hfe00;
			16'h9a62: y = 16'hfe00;
			16'h9a63: y = 16'hfe00;
			16'h9a64: y = 16'hfe00;
			16'h9a65: y = 16'hfe00;
			16'h9a66: y = 16'hfe00;
			16'h9a67: y = 16'hfe00;
			16'h9a68: y = 16'hfe00;
			16'h9a69: y = 16'hfe00;
			16'h9a6a: y = 16'hfe00;
			16'h9a6b: y = 16'hfe00;
			16'h9a6c: y = 16'hfe00;
			16'h9a6d: y = 16'hfe00;
			16'h9a6e: y = 16'hfe00;
			16'h9a6f: y = 16'hfe00;
			16'h9a70: y = 16'hfe00;
			16'h9a71: y = 16'hfe00;
			16'h9a72: y = 16'hfe00;
			16'h9a73: y = 16'hfe00;
			16'h9a74: y = 16'hfe00;
			16'h9a75: y = 16'hfe00;
			16'h9a76: y = 16'hfe00;
			16'h9a77: y = 16'hfe00;
			16'h9a78: y = 16'hfe00;
			16'h9a79: y = 16'hfe00;
			16'h9a7a: y = 16'hfe00;
			16'h9a7b: y = 16'hfe00;
			16'h9a7c: y = 16'hfe00;
			16'h9a7d: y = 16'hfe00;
			16'h9a7e: y = 16'hfe00;
			16'h9a7f: y = 16'hfe00;
			16'h9a80: y = 16'hfe00;
			16'h9a81: y = 16'hfe00;
			16'h9a82: y = 16'hfe00;
			16'h9a83: y = 16'hfe00;
			16'h9a84: y = 16'hfe00;
			16'h9a85: y = 16'hfe00;
			16'h9a86: y = 16'hfe00;
			16'h9a87: y = 16'hfe00;
			16'h9a88: y = 16'hfe00;
			16'h9a89: y = 16'hfe00;
			16'h9a8a: y = 16'hfe00;
			16'h9a8b: y = 16'hfe00;
			16'h9a8c: y = 16'hfe00;
			16'h9a8d: y = 16'hfe00;
			16'h9a8e: y = 16'hfe00;
			16'h9a8f: y = 16'hfe00;
			16'h9a90: y = 16'hfe00;
			16'h9a91: y = 16'hfe00;
			16'h9a92: y = 16'hfe00;
			16'h9a93: y = 16'hfe00;
			16'h9a94: y = 16'hfe00;
			16'h9a95: y = 16'hfe00;
			16'h9a96: y = 16'hfe00;
			16'h9a97: y = 16'hfe00;
			16'h9a98: y = 16'hfe00;
			16'h9a99: y = 16'hfe00;
			16'h9a9a: y = 16'hfe00;
			16'h9a9b: y = 16'hfe00;
			16'h9a9c: y = 16'hfe00;
			16'h9a9d: y = 16'hfe00;
			16'h9a9e: y = 16'hfe00;
			16'h9a9f: y = 16'hfe00;
			16'h9aa0: y = 16'hfe00;
			16'h9aa1: y = 16'hfe00;
			16'h9aa2: y = 16'hfe00;
			16'h9aa3: y = 16'hfe00;
			16'h9aa4: y = 16'hfe00;
			16'h9aa5: y = 16'hfe00;
			16'h9aa6: y = 16'hfe00;
			16'h9aa7: y = 16'hfe00;
			16'h9aa8: y = 16'hfe00;
			16'h9aa9: y = 16'hfe00;
			16'h9aaa: y = 16'hfe00;
			16'h9aab: y = 16'hfe00;
			16'h9aac: y = 16'hfe00;
			16'h9aad: y = 16'hfe00;
			16'h9aae: y = 16'hfe00;
			16'h9aaf: y = 16'hfe00;
			16'h9ab0: y = 16'hfe00;
			16'h9ab1: y = 16'hfe00;
			16'h9ab2: y = 16'hfe00;
			16'h9ab3: y = 16'hfe00;
			16'h9ab4: y = 16'hfe00;
			16'h9ab5: y = 16'hfe00;
			16'h9ab6: y = 16'hfe00;
			16'h9ab7: y = 16'hfe00;
			16'h9ab8: y = 16'hfe00;
			16'h9ab9: y = 16'hfe00;
			16'h9aba: y = 16'hfe00;
			16'h9abb: y = 16'hfe00;
			16'h9abc: y = 16'hfe00;
			16'h9abd: y = 16'hfe00;
			16'h9abe: y = 16'hfe00;
			16'h9abf: y = 16'hfe00;
			16'h9ac0: y = 16'hfe00;
			16'h9ac1: y = 16'hfe00;
			16'h9ac2: y = 16'hfe00;
			16'h9ac3: y = 16'hfe00;
			16'h9ac4: y = 16'hfe00;
			16'h9ac5: y = 16'hfe00;
			16'h9ac6: y = 16'hfe00;
			16'h9ac7: y = 16'hfe00;
			16'h9ac8: y = 16'hfe00;
			16'h9ac9: y = 16'hfe00;
			16'h9aca: y = 16'hfe00;
			16'h9acb: y = 16'hfe00;
			16'h9acc: y = 16'hfe00;
			16'h9acd: y = 16'hfe00;
			16'h9ace: y = 16'hfe00;
			16'h9acf: y = 16'hfe00;
			16'h9ad0: y = 16'hfe00;
			16'h9ad1: y = 16'hfe00;
			16'h9ad2: y = 16'hfe00;
			16'h9ad3: y = 16'hfe00;
			16'h9ad4: y = 16'hfe00;
			16'h9ad5: y = 16'hfe00;
			16'h9ad6: y = 16'hfe00;
			16'h9ad7: y = 16'hfe00;
			16'h9ad8: y = 16'hfe00;
			16'h9ad9: y = 16'hfe00;
			16'h9ada: y = 16'hfe00;
			16'h9adb: y = 16'hfe00;
			16'h9adc: y = 16'hfe00;
			16'h9add: y = 16'hfe00;
			16'h9ade: y = 16'hfe00;
			16'h9adf: y = 16'hfe00;
			16'h9ae0: y = 16'hfe00;
			16'h9ae1: y = 16'hfe00;
			16'h9ae2: y = 16'hfe00;
			16'h9ae3: y = 16'hfe00;
			16'h9ae4: y = 16'hfe00;
			16'h9ae5: y = 16'hfe00;
			16'h9ae6: y = 16'hfe00;
			16'h9ae7: y = 16'hfe00;
			16'h9ae8: y = 16'hfe00;
			16'h9ae9: y = 16'hfe00;
			16'h9aea: y = 16'hfe00;
			16'h9aeb: y = 16'hfe00;
			16'h9aec: y = 16'hfe00;
			16'h9aed: y = 16'hfe00;
			16'h9aee: y = 16'hfe00;
			16'h9aef: y = 16'hfe00;
			16'h9af0: y = 16'hfe00;
			16'h9af1: y = 16'hfe00;
			16'h9af2: y = 16'hfe00;
			16'h9af3: y = 16'hfe00;
			16'h9af4: y = 16'hfe00;
			16'h9af5: y = 16'hfe00;
			16'h9af6: y = 16'hfe00;
			16'h9af7: y = 16'hfe00;
			16'h9af8: y = 16'hfe00;
			16'h9af9: y = 16'hfe00;
			16'h9afa: y = 16'hfe00;
			16'h9afb: y = 16'hfe00;
			16'h9afc: y = 16'hfe00;
			16'h9afd: y = 16'hfe00;
			16'h9afe: y = 16'hfe00;
			16'h9aff: y = 16'hfe00;
			16'h9b00: y = 16'hfe00;
			16'h9b01: y = 16'hfe00;
			16'h9b02: y = 16'hfe00;
			16'h9b03: y = 16'hfe00;
			16'h9b04: y = 16'hfe00;
			16'h9b05: y = 16'hfe00;
			16'h9b06: y = 16'hfe00;
			16'h9b07: y = 16'hfe00;
			16'h9b08: y = 16'hfe00;
			16'h9b09: y = 16'hfe00;
			16'h9b0a: y = 16'hfe00;
			16'h9b0b: y = 16'hfe00;
			16'h9b0c: y = 16'hfe00;
			16'h9b0d: y = 16'hfe00;
			16'h9b0e: y = 16'hfe00;
			16'h9b0f: y = 16'hfe00;
			16'h9b10: y = 16'hfe00;
			16'h9b11: y = 16'hfe00;
			16'h9b12: y = 16'hfe00;
			16'h9b13: y = 16'hfe00;
			16'h9b14: y = 16'hfe00;
			16'h9b15: y = 16'hfe00;
			16'h9b16: y = 16'hfe00;
			16'h9b17: y = 16'hfe00;
			16'h9b18: y = 16'hfe00;
			16'h9b19: y = 16'hfe00;
			16'h9b1a: y = 16'hfe00;
			16'h9b1b: y = 16'hfe00;
			16'h9b1c: y = 16'hfe00;
			16'h9b1d: y = 16'hfe00;
			16'h9b1e: y = 16'hfe00;
			16'h9b1f: y = 16'hfe00;
			16'h9b20: y = 16'hfe00;
			16'h9b21: y = 16'hfe00;
			16'h9b22: y = 16'hfe00;
			16'h9b23: y = 16'hfe00;
			16'h9b24: y = 16'hfe00;
			16'h9b25: y = 16'hfe00;
			16'h9b26: y = 16'hfe00;
			16'h9b27: y = 16'hfe00;
			16'h9b28: y = 16'hfe00;
			16'h9b29: y = 16'hfe00;
			16'h9b2a: y = 16'hfe00;
			16'h9b2b: y = 16'hfe00;
			16'h9b2c: y = 16'hfe00;
			16'h9b2d: y = 16'hfe00;
			16'h9b2e: y = 16'hfe00;
			16'h9b2f: y = 16'hfe00;
			16'h9b30: y = 16'hfe00;
			16'h9b31: y = 16'hfe00;
			16'h9b32: y = 16'hfe00;
			16'h9b33: y = 16'hfe00;
			16'h9b34: y = 16'hfe00;
			16'h9b35: y = 16'hfe00;
			16'h9b36: y = 16'hfe00;
			16'h9b37: y = 16'hfe00;
			16'h9b38: y = 16'hfe00;
			16'h9b39: y = 16'hfe00;
			16'h9b3a: y = 16'hfe00;
			16'h9b3b: y = 16'hfe00;
			16'h9b3c: y = 16'hfe00;
			16'h9b3d: y = 16'hfe00;
			16'h9b3e: y = 16'hfe00;
			16'h9b3f: y = 16'hfe00;
			16'h9b40: y = 16'hfe00;
			16'h9b41: y = 16'hfe00;
			16'h9b42: y = 16'hfe00;
			16'h9b43: y = 16'hfe00;
			16'h9b44: y = 16'hfe00;
			16'h9b45: y = 16'hfe00;
			16'h9b46: y = 16'hfe00;
			16'h9b47: y = 16'hfe00;
			16'h9b48: y = 16'hfe00;
			16'h9b49: y = 16'hfe00;
			16'h9b4a: y = 16'hfe00;
			16'h9b4b: y = 16'hfe00;
			16'h9b4c: y = 16'hfe00;
			16'h9b4d: y = 16'hfe00;
			16'h9b4e: y = 16'hfe00;
			16'h9b4f: y = 16'hfe00;
			16'h9b50: y = 16'hfe00;
			16'h9b51: y = 16'hfe00;
			16'h9b52: y = 16'hfe00;
			16'h9b53: y = 16'hfe00;
			16'h9b54: y = 16'hfe00;
			16'h9b55: y = 16'hfe00;
			16'h9b56: y = 16'hfe00;
			16'h9b57: y = 16'hfe00;
			16'h9b58: y = 16'hfe00;
			16'h9b59: y = 16'hfe00;
			16'h9b5a: y = 16'hfe00;
			16'h9b5b: y = 16'hfe00;
			16'h9b5c: y = 16'hfe00;
			16'h9b5d: y = 16'hfe00;
			16'h9b5e: y = 16'hfe00;
			16'h9b5f: y = 16'hfe00;
			16'h9b60: y = 16'hfe00;
			16'h9b61: y = 16'hfe00;
			16'h9b62: y = 16'hfe00;
			16'h9b63: y = 16'hfe00;
			16'h9b64: y = 16'hfe00;
			16'h9b65: y = 16'hfe00;
			16'h9b66: y = 16'hfe00;
			16'h9b67: y = 16'hfe00;
			16'h9b68: y = 16'hfe00;
			16'h9b69: y = 16'hfe00;
			16'h9b6a: y = 16'hfe00;
			16'h9b6b: y = 16'hfe00;
			16'h9b6c: y = 16'hfe00;
			16'h9b6d: y = 16'hfe00;
			16'h9b6e: y = 16'hfe00;
			16'h9b6f: y = 16'hfe00;
			16'h9b70: y = 16'hfe00;
			16'h9b71: y = 16'hfe00;
			16'h9b72: y = 16'hfe00;
			16'h9b73: y = 16'hfe00;
			16'h9b74: y = 16'hfe00;
			16'h9b75: y = 16'hfe00;
			16'h9b76: y = 16'hfe00;
			16'h9b77: y = 16'hfe00;
			16'h9b78: y = 16'hfe00;
			16'h9b79: y = 16'hfe00;
			16'h9b7a: y = 16'hfe00;
			16'h9b7b: y = 16'hfe00;
			16'h9b7c: y = 16'hfe00;
			16'h9b7d: y = 16'hfe00;
			16'h9b7e: y = 16'hfe00;
			16'h9b7f: y = 16'hfe00;
			16'h9b80: y = 16'hfe00;
			16'h9b81: y = 16'hfe00;
			16'h9b82: y = 16'hfe00;
			16'h9b83: y = 16'hfe00;
			16'h9b84: y = 16'hfe00;
			16'h9b85: y = 16'hfe00;
			16'h9b86: y = 16'hfe00;
			16'h9b87: y = 16'hfe00;
			16'h9b88: y = 16'hfe00;
			16'h9b89: y = 16'hfe00;
			16'h9b8a: y = 16'hfe00;
			16'h9b8b: y = 16'hfe00;
			16'h9b8c: y = 16'hfe00;
			16'h9b8d: y = 16'hfe00;
			16'h9b8e: y = 16'hfe00;
			16'h9b8f: y = 16'hfe00;
			16'h9b90: y = 16'hfe00;
			16'h9b91: y = 16'hfe00;
			16'h9b92: y = 16'hfe00;
			16'h9b93: y = 16'hfe00;
			16'h9b94: y = 16'hfe00;
			16'h9b95: y = 16'hfe00;
			16'h9b96: y = 16'hfe00;
			16'h9b97: y = 16'hfe00;
			16'h9b98: y = 16'hfe00;
			16'h9b99: y = 16'hfe00;
			16'h9b9a: y = 16'hfe00;
			16'h9b9b: y = 16'hfe00;
			16'h9b9c: y = 16'hfe00;
			16'h9b9d: y = 16'hfe00;
			16'h9b9e: y = 16'hfe00;
			16'h9b9f: y = 16'hfe00;
			16'h9ba0: y = 16'hfe00;
			16'h9ba1: y = 16'hfe00;
			16'h9ba2: y = 16'hfe00;
			16'h9ba3: y = 16'hfe00;
			16'h9ba4: y = 16'hfe00;
			16'h9ba5: y = 16'hfe00;
			16'h9ba6: y = 16'hfe00;
			16'h9ba7: y = 16'hfe00;
			16'h9ba8: y = 16'hfe00;
			16'h9ba9: y = 16'hfe00;
			16'h9baa: y = 16'hfe00;
			16'h9bab: y = 16'hfe00;
			16'h9bac: y = 16'hfe00;
			16'h9bad: y = 16'hfe00;
			16'h9bae: y = 16'hfe00;
			16'h9baf: y = 16'hfe00;
			16'h9bb0: y = 16'hfe00;
			16'h9bb1: y = 16'hfe00;
			16'h9bb2: y = 16'hfe00;
			16'h9bb3: y = 16'hfe00;
			16'h9bb4: y = 16'hfe00;
			16'h9bb5: y = 16'hfe00;
			16'h9bb6: y = 16'hfe00;
			16'h9bb7: y = 16'hfe00;
			16'h9bb8: y = 16'hfe00;
			16'h9bb9: y = 16'hfe00;
			16'h9bba: y = 16'hfe00;
			16'h9bbb: y = 16'hfe00;
			16'h9bbc: y = 16'hfe00;
			16'h9bbd: y = 16'hfe00;
			16'h9bbe: y = 16'hfe00;
			16'h9bbf: y = 16'hfe00;
			16'h9bc0: y = 16'hfe00;
			16'h9bc1: y = 16'hfe00;
			16'h9bc2: y = 16'hfe00;
			16'h9bc3: y = 16'hfe00;
			16'h9bc4: y = 16'hfe00;
			16'h9bc5: y = 16'hfe00;
			16'h9bc6: y = 16'hfe00;
			16'h9bc7: y = 16'hfe00;
			16'h9bc8: y = 16'hfe00;
			16'h9bc9: y = 16'hfe00;
			16'h9bca: y = 16'hfe00;
			16'h9bcb: y = 16'hfe00;
			16'h9bcc: y = 16'hfe00;
			16'h9bcd: y = 16'hfe00;
			16'h9bce: y = 16'hfe00;
			16'h9bcf: y = 16'hfe00;
			16'h9bd0: y = 16'hfe00;
			16'h9bd1: y = 16'hfe00;
			16'h9bd2: y = 16'hfe00;
			16'h9bd3: y = 16'hfe00;
			16'h9bd4: y = 16'hfe00;
			16'h9bd5: y = 16'hfe00;
			16'h9bd6: y = 16'hfe00;
			16'h9bd7: y = 16'hfe00;
			16'h9bd8: y = 16'hfe00;
			16'h9bd9: y = 16'hfe00;
			16'h9bda: y = 16'hfe00;
			16'h9bdb: y = 16'hfe00;
			16'h9bdc: y = 16'hfe00;
			16'h9bdd: y = 16'hfe00;
			16'h9bde: y = 16'hfe00;
			16'h9bdf: y = 16'hfe00;
			16'h9be0: y = 16'hfe00;
			16'h9be1: y = 16'hfe00;
			16'h9be2: y = 16'hfe00;
			16'h9be3: y = 16'hfe00;
			16'h9be4: y = 16'hfe00;
			16'h9be5: y = 16'hfe00;
			16'h9be6: y = 16'hfe00;
			16'h9be7: y = 16'hfe00;
			16'h9be8: y = 16'hfe00;
			16'h9be9: y = 16'hfe00;
			16'h9bea: y = 16'hfe00;
			16'h9beb: y = 16'hfe00;
			16'h9bec: y = 16'hfe00;
			16'h9bed: y = 16'hfe00;
			16'h9bee: y = 16'hfe00;
			16'h9bef: y = 16'hfe00;
			16'h9bf0: y = 16'hfe00;
			16'h9bf1: y = 16'hfe00;
			16'h9bf2: y = 16'hfe00;
			16'h9bf3: y = 16'hfe00;
			16'h9bf4: y = 16'hfe00;
			16'h9bf5: y = 16'hfe00;
			16'h9bf6: y = 16'hfe00;
			16'h9bf7: y = 16'hfe00;
			16'h9bf8: y = 16'hfe00;
			16'h9bf9: y = 16'hfe00;
			16'h9bfa: y = 16'hfe00;
			16'h9bfb: y = 16'hfe00;
			16'h9bfc: y = 16'hfe00;
			16'h9bfd: y = 16'hfe00;
			16'h9bfe: y = 16'hfe00;
			16'h9bff: y = 16'hfe00;
			16'h9c00: y = 16'hfe00;
			16'h9c01: y = 16'hfe00;
			16'h9c02: y = 16'hfe00;
			16'h9c03: y = 16'hfe00;
			16'h9c04: y = 16'hfe00;
			16'h9c05: y = 16'hfe00;
			16'h9c06: y = 16'hfe00;
			16'h9c07: y = 16'hfe00;
			16'h9c08: y = 16'hfe00;
			16'h9c09: y = 16'hfe00;
			16'h9c0a: y = 16'hfe00;
			16'h9c0b: y = 16'hfe00;
			16'h9c0c: y = 16'hfe00;
			16'h9c0d: y = 16'hfe00;
			16'h9c0e: y = 16'hfe00;
			16'h9c0f: y = 16'hfe00;
			16'h9c10: y = 16'hfe00;
			16'h9c11: y = 16'hfe00;
			16'h9c12: y = 16'hfe00;
			16'h9c13: y = 16'hfe00;
			16'h9c14: y = 16'hfe00;
			16'h9c15: y = 16'hfe00;
			16'h9c16: y = 16'hfe00;
			16'h9c17: y = 16'hfe00;
			16'h9c18: y = 16'hfe00;
			16'h9c19: y = 16'hfe00;
			16'h9c1a: y = 16'hfe00;
			16'h9c1b: y = 16'hfe00;
			16'h9c1c: y = 16'hfe00;
			16'h9c1d: y = 16'hfe00;
			16'h9c1e: y = 16'hfe00;
			16'h9c1f: y = 16'hfe00;
			16'h9c20: y = 16'hfe00;
			16'h9c21: y = 16'hfe00;
			16'h9c22: y = 16'hfe00;
			16'h9c23: y = 16'hfe00;
			16'h9c24: y = 16'hfe00;
			16'h9c25: y = 16'hfe00;
			16'h9c26: y = 16'hfe00;
			16'h9c27: y = 16'hfe00;
			16'h9c28: y = 16'hfe00;
			16'h9c29: y = 16'hfe00;
			16'h9c2a: y = 16'hfe00;
			16'h9c2b: y = 16'hfe00;
			16'h9c2c: y = 16'hfe00;
			16'h9c2d: y = 16'hfe00;
			16'h9c2e: y = 16'hfe00;
			16'h9c2f: y = 16'hfe00;
			16'h9c30: y = 16'hfe00;
			16'h9c31: y = 16'hfe00;
			16'h9c32: y = 16'hfe00;
			16'h9c33: y = 16'hfe00;
			16'h9c34: y = 16'hfe00;
			16'h9c35: y = 16'hfe00;
			16'h9c36: y = 16'hfe00;
			16'h9c37: y = 16'hfe00;
			16'h9c38: y = 16'hfe00;
			16'h9c39: y = 16'hfe00;
			16'h9c3a: y = 16'hfe00;
			16'h9c3b: y = 16'hfe00;
			16'h9c3c: y = 16'hfe00;
			16'h9c3d: y = 16'hfe00;
			16'h9c3e: y = 16'hfe00;
			16'h9c3f: y = 16'hfe00;
			16'h9c40: y = 16'hfe00;
			16'h9c41: y = 16'hfe00;
			16'h9c42: y = 16'hfe00;
			16'h9c43: y = 16'hfe00;
			16'h9c44: y = 16'hfe00;
			16'h9c45: y = 16'hfe00;
			16'h9c46: y = 16'hfe00;
			16'h9c47: y = 16'hfe00;
			16'h9c48: y = 16'hfe00;
			16'h9c49: y = 16'hfe00;
			16'h9c4a: y = 16'hfe00;
			16'h9c4b: y = 16'hfe00;
			16'h9c4c: y = 16'hfe00;
			16'h9c4d: y = 16'hfe00;
			16'h9c4e: y = 16'hfe00;
			16'h9c4f: y = 16'hfe00;
			16'h9c50: y = 16'hfe00;
			16'h9c51: y = 16'hfe00;
			16'h9c52: y = 16'hfe00;
			16'h9c53: y = 16'hfe00;
			16'h9c54: y = 16'hfe00;
			16'h9c55: y = 16'hfe00;
			16'h9c56: y = 16'hfe00;
			16'h9c57: y = 16'hfe00;
			16'h9c58: y = 16'hfe00;
			16'h9c59: y = 16'hfe00;
			16'h9c5a: y = 16'hfe00;
			16'h9c5b: y = 16'hfe00;
			16'h9c5c: y = 16'hfe00;
			16'h9c5d: y = 16'hfe00;
			16'h9c5e: y = 16'hfe00;
			16'h9c5f: y = 16'hfe00;
			16'h9c60: y = 16'hfe00;
			16'h9c61: y = 16'hfe00;
			16'h9c62: y = 16'hfe00;
			16'h9c63: y = 16'hfe00;
			16'h9c64: y = 16'hfe00;
			16'h9c65: y = 16'hfe00;
			16'h9c66: y = 16'hfe00;
			16'h9c67: y = 16'hfe00;
			16'h9c68: y = 16'hfe00;
			16'h9c69: y = 16'hfe00;
			16'h9c6a: y = 16'hfe00;
			16'h9c6b: y = 16'hfe00;
			16'h9c6c: y = 16'hfe00;
			16'h9c6d: y = 16'hfe00;
			16'h9c6e: y = 16'hfe00;
			16'h9c6f: y = 16'hfe00;
			16'h9c70: y = 16'hfe00;
			16'h9c71: y = 16'hfe00;
			16'h9c72: y = 16'hfe00;
			16'h9c73: y = 16'hfe00;
			16'h9c74: y = 16'hfe00;
			16'h9c75: y = 16'hfe00;
			16'h9c76: y = 16'hfe00;
			16'h9c77: y = 16'hfe00;
			16'h9c78: y = 16'hfe00;
			16'h9c79: y = 16'hfe00;
			16'h9c7a: y = 16'hfe00;
			16'h9c7b: y = 16'hfe00;
			16'h9c7c: y = 16'hfe00;
			16'h9c7d: y = 16'hfe00;
			16'h9c7e: y = 16'hfe00;
			16'h9c7f: y = 16'hfe00;
			16'h9c80: y = 16'hfe00;
			16'h9c81: y = 16'hfe00;
			16'h9c82: y = 16'hfe00;
			16'h9c83: y = 16'hfe00;
			16'h9c84: y = 16'hfe00;
			16'h9c85: y = 16'hfe00;
			16'h9c86: y = 16'hfe00;
			16'h9c87: y = 16'hfe00;
			16'h9c88: y = 16'hfe00;
			16'h9c89: y = 16'hfe00;
			16'h9c8a: y = 16'hfe00;
			16'h9c8b: y = 16'hfe00;
			16'h9c8c: y = 16'hfe00;
			16'h9c8d: y = 16'hfe00;
			16'h9c8e: y = 16'hfe00;
			16'h9c8f: y = 16'hfe00;
			16'h9c90: y = 16'hfe00;
			16'h9c91: y = 16'hfe00;
			16'h9c92: y = 16'hfe00;
			16'h9c93: y = 16'hfe00;
			16'h9c94: y = 16'hfe00;
			16'h9c95: y = 16'hfe00;
			16'h9c96: y = 16'hfe00;
			16'h9c97: y = 16'hfe00;
			16'h9c98: y = 16'hfe00;
			16'h9c99: y = 16'hfe00;
			16'h9c9a: y = 16'hfe00;
			16'h9c9b: y = 16'hfe00;
			16'h9c9c: y = 16'hfe00;
			16'h9c9d: y = 16'hfe00;
			16'h9c9e: y = 16'hfe00;
			16'h9c9f: y = 16'hfe00;
			16'h9ca0: y = 16'hfe00;
			16'h9ca1: y = 16'hfe00;
			16'h9ca2: y = 16'hfe00;
			16'h9ca3: y = 16'hfe00;
			16'h9ca4: y = 16'hfe00;
			16'h9ca5: y = 16'hfe00;
			16'h9ca6: y = 16'hfe00;
			16'h9ca7: y = 16'hfe00;
			16'h9ca8: y = 16'hfe00;
			16'h9ca9: y = 16'hfe00;
			16'h9caa: y = 16'hfe00;
			16'h9cab: y = 16'hfe00;
			16'h9cac: y = 16'hfe00;
			16'h9cad: y = 16'hfe00;
			16'h9cae: y = 16'hfe00;
			16'h9caf: y = 16'hfe00;
			16'h9cb0: y = 16'hfe00;
			16'h9cb1: y = 16'hfe00;
			16'h9cb2: y = 16'hfe00;
			16'h9cb3: y = 16'hfe00;
			16'h9cb4: y = 16'hfe00;
			16'h9cb5: y = 16'hfe00;
			16'h9cb6: y = 16'hfe00;
			16'h9cb7: y = 16'hfe00;
			16'h9cb8: y = 16'hfe00;
			16'h9cb9: y = 16'hfe00;
			16'h9cba: y = 16'hfe00;
			16'h9cbb: y = 16'hfe00;
			16'h9cbc: y = 16'hfe00;
			16'h9cbd: y = 16'hfe00;
			16'h9cbe: y = 16'hfe00;
			16'h9cbf: y = 16'hfe00;
			16'h9cc0: y = 16'hfe00;
			16'h9cc1: y = 16'hfe00;
			16'h9cc2: y = 16'hfe00;
			16'h9cc3: y = 16'hfe00;
			16'h9cc4: y = 16'hfe00;
			16'h9cc5: y = 16'hfe00;
			16'h9cc6: y = 16'hfe00;
			16'h9cc7: y = 16'hfe00;
			16'h9cc8: y = 16'hfe00;
			16'h9cc9: y = 16'hfe00;
			16'h9cca: y = 16'hfe00;
			16'h9ccb: y = 16'hfe00;
			16'h9ccc: y = 16'hfe00;
			16'h9ccd: y = 16'hfe00;
			16'h9cce: y = 16'hfe00;
			16'h9ccf: y = 16'hfe00;
			16'h9cd0: y = 16'hfe00;
			16'h9cd1: y = 16'hfe00;
			16'h9cd2: y = 16'hfe00;
			16'h9cd3: y = 16'hfe00;
			16'h9cd4: y = 16'hfe00;
			16'h9cd5: y = 16'hfe00;
			16'h9cd6: y = 16'hfe00;
			16'h9cd7: y = 16'hfe00;
			16'h9cd8: y = 16'hfe00;
			16'h9cd9: y = 16'hfe00;
			16'h9cda: y = 16'hfe00;
			16'h9cdb: y = 16'hfe00;
			16'h9cdc: y = 16'hfe00;
			16'h9cdd: y = 16'hfe00;
			16'h9cde: y = 16'hfe00;
			16'h9cdf: y = 16'hfe00;
			16'h9ce0: y = 16'hfe00;
			16'h9ce1: y = 16'hfe00;
			16'h9ce2: y = 16'hfe00;
			16'h9ce3: y = 16'hfe00;
			16'h9ce4: y = 16'hfe00;
			16'h9ce5: y = 16'hfe00;
			16'h9ce6: y = 16'hfe00;
			16'h9ce7: y = 16'hfe00;
			16'h9ce8: y = 16'hfe00;
			16'h9ce9: y = 16'hfe00;
			16'h9cea: y = 16'hfe00;
			16'h9ceb: y = 16'hfe00;
			16'h9cec: y = 16'hfe00;
			16'h9ced: y = 16'hfe00;
			16'h9cee: y = 16'hfe00;
			16'h9cef: y = 16'hfe00;
			16'h9cf0: y = 16'hfe00;
			16'h9cf1: y = 16'hfe00;
			16'h9cf2: y = 16'hfe00;
			16'h9cf3: y = 16'hfe00;
			16'h9cf4: y = 16'hfe00;
			16'h9cf5: y = 16'hfe00;
			16'h9cf6: y = 16'hfe00;
			16'h9cf7: y = 16'hfe00;
			16'h9cf8: y = 16'hfe00;
			16'h9cf9: y = 16'hfe00;
			16'h9cfa: y = 16'hfe00;
			16'h9cfb: y = 16'hfe00;
			16'h9cfc: y = 16'hfe00;
			16'h9cfd: y = 16'hfe00;
			16'h9cfe: y = 16'hfe00;
			16'h9cff: y = 16'hfe00;
			16'h9d00: y = 16'hfe00;
			16'h9d01: y = 16'hfe00;
			16'h9d02: y = 16'hfe00;
			16'h9d03: y = 16'hfe00;
			16'h9d04: y = 16'hfe00;
			16'h9d05: y = 16'hfe00;
			16'h9d06: y = 16'hfe00;
			16'h9d07: y = 16'hfe00;
			16'h9d08: y = 16'hfe00;
			16'h9d09: y = 16'hfe00;
			16'h9d0a: y = 16'hfe00;
			16'h9d0b: y = 16'hfe00;
			16'h9d0c: y = 16'hfe00;
			16'h9d0d: y = 16'hfe00;
			16'h9d0e: y = 16'hfe00;
			16'h9d0f: y = 16'hfe00;
			16'h9d10: y = 16'hfe00;
			16'h9d11: y = 16'hfe00;
			16'h9d12: y = 16'hfe00;
			16'h9d13: y = 16'hfe00;
			16'h9d14: y = 16'hfe00;
			16'h9d15: y = 16'hfe00;
			16'h9d16: y = 16'hfe00;
			16'h9d17: y = 16'hfe00;
			16'h9d18: y = 16'hfe00;
			16'h9d19: y = 16'hfe00;
			16'h9d1a: y = 16'hfe00;
			16'h9d1b: y = 16'hfe00;
			16'h9d1c: y = 16'hfe00;
			16'h9d1d: y = 16'hfe00;
			16'h9d1e: y = 16'hfe00;
			16'h9d1f: y = 16'hfe00;
			16'h9d20: y = 16'hfe00;
			16'h9d21: y = 16'hfe00;
			16'h9d22: y = 16'hfe00;
			16'h9d23: y = 16'hfe00;
			16'h9d24: y = 16'hfe00;
			16'h9d25: y = 16'hfe00;
			16'h9d26: y = 16'hfe00;
			16'h9d27: y = 16'hfe00;
			16'h9d28: y = 16'hfe00;
			16'h9d29: y = 16'hfe00;
			16'h9d2a: y = 16'hfe00;
			16'h9d2b: y = 16'hfe00;
			16'h9d2c: y = 16'hfe00;
			16'h9d2d: y = 16'hfe00;
			16'h9d2e: y = 16'hfe00;
			16'h9d2f: y = 16'hfe00;
			16'h9d30: y = 16'hfe00;
			16'h9d31: y = 16'hfe00;
			16'h9d32: y = 16'hfe00;
			16'h9d33: y = 16'hfe00;
			16'h9d34: y = 16'hfe00;
			16'h9d35: y = 16'hfe00;
			16'h9d36: y = 16'hfe00;
			16'h9d37: y = 16'hfe00;
			16'h9d38: y = 16'hfe00;
			16'h9d39: y = 16'hfe00;
			16'h9d3a: y = 16'hfe00;
			16'h9d3b: y = 16'hfe00;
			16'h9d3c: y = 16'hfe00;
			16'h9d3d: y = 16'hfe00;
			16'h9d3e: y = 16'hfe00;
			16'h9d3f: y = 16'hfe00;
			16'h9d40: y = 16'hfe00;
			16'h9d41: y = 16'hfe00;
			16'h9d42: y = 16'hfe00;
			16'h9d43: y = 16'hfe00;
			16'h9d44: y = 16'hfe00;
			16'h9d45: y = 16'hfe00;
			16'h9d46: y = 16'hfe00;
			16'h9d47: y = 16'hfe00;
			16'h9d48: y = 16'hfe00;
			16'h9d49: y = 16'hfe00;
			16'h9d4a: y = 16'hfe00;
			16'h9d4b: y = 16'hfe00;
			16'h9d4c: y = 16'hfe00;
			16'h9d4d: y = 16'hfe00;
			16'h9d4e: y = 16'hfe00;
			16'h9d4f: y = 16'hfe00;
			16'h9d50: y = 16'hfe00;
			16'h9d51: y = 16'hfe00;
			16'h9d52: y = 16'hfe00;
			16'h9d53: y = 16'hfe00;
			16'h9d54: y = 16'hfe00;
			16'h9d55: y = 16'hfe00;
			16'h9d56: y = 16'hfe00;
			16'h9d57: y = 16'hfe00;
			16'h9d58: y = 16'hfe00;
			16'h9d59: y = 16'hfe00;
			16'h9d5a: y = 16'hfe00;
			16'h9d5b: y = 16'hfe00;
			16'h9d5c: y = 16'hfe00;
			16'h9d5d: y = 16'hfe00;
			16'h9d5e: y = 16'hfe00;
			16'h9d5f: y = 16'hfe00;
			16'h9d60: y = 16'hfe00;
			16'h9d61: y = 16'hfe00;
			16'h9d62: y = 16'hfe00;
			16'h9d63: y = 16'hfe00;
			16'h9d64: y = 16'hfe00;
			16'h9d65: y = 16'hfe00;
			16'h9d66: y = 16'hfe00;
			16'h9d67: y = 16'hfe00;
			16'h9d68: y = 16'hfe00;
			16'h9d69: y = 16'hfe00;
			16'h9d6a: y = 16'hfe00;
			16'h9d6b: y = 16'hfe00;
			16'h9d6c: y = 16'hfe00;
			16'h9d6d: y = 16'hfe00;
			16'h9d6e: y = 16'hfe00;
			16'h9d6f: y = 16'hfe00;
			16'h9d70: y = 16'hfe00;
			16'h9d71: y = 16'hfe00;
			16'h9d72: y = 16'hfe00;
			16'h9d73: y = 16'hfe00;
			16'h9d74: y = 16'hfe00;
			16'h9d75: y = 16'hfe00;
			16'h9d76: y = 16'hfe00;
			16'h9d77: y = 16'hfe00;
			16'h9d78: y = 16'hfe00;
			16'h9d79: y = 16'hfe00;
			16'h9d7a: y = 16'hfe00;
			16'h9d7b: y = 16'hfe00;
			16'h9d7c: y = 16'hfe00;
			16'h9d7d: y = 16'hfe00;
			16'h9d7e: y = 16'hfe00;
			16'h9d7f: y = 16'hfe00;
			16'h9d80: y = 16'hfe00;
			16'h9d81: y = 16'hfe00;
			16'h9d82: y = 16'hfe00;
			16'h9d83: y = 16'hfe00;
			16'h9d84: y = 16'hfe00;
			16'h9d85: y = 16'hfe00;
			16'h9d86: y = 16'hfe00;
			16'h9d87: y = 16'hfe00;
			16'h9d88: y = 16'hfe00;
			16'h9d89: y = 16'hfe00;
			16'h9d8a: y = 16'hfe00;
			16'h9d8b: y = 16'hfe00;
			16'h9d8c: y = 16'hfe00;
			16'h9d8d: y = 16'hfe00;
			16'h9d8e: y = 16'hfe00;
			16'h9d8f: y = 16'hfe00;
			16'h9d90: y = 16'hfe00;
			16'h9d91: y = 16'hfe00;
			16'h9d92: y = 16'hfe00;
			16'h9d93: y = 16'hfe00;
			16'h9d94: y = 16'hfe00;
			16'h9d95: y = 16'hfe00;
			16'h9d96: y = 16'hfe00;
			16'h9d97: y = 16'hfe00;
			16'h9d98: y = 16'hfe00;
			16'h9d99: y = 16'hfe00;
			16'h9d9a: y = 16'hfe00;
			16'h9d9b: y = 16'hfe00;
			16'h9d9c: y = 16'hfe00;
			16'h9d9d: y = 16'hfe00;
			16'h9d9e: y = 16'hfe00;
			16'h9d9f: y = 16'hfe00;
			16'h9da0: y = 16'hfe00;
			16'h9da1: y = 16'hfe00;
			16'h9da2: y = 16'hfe00;
			16'h9da3: y = 16'hfe00;
			16'h9da4: y = 16'hfe00;
			16'h9da5: y = 16'hfe00;
			16'h9da6: y = 16'hfe00;
			16'h9da7: y = 16'hfe00;
			16'h9da8: y = 16'hfe00;
			16'h9da9: y = 16'hfe00;
			16'h9daa: y = 16'hfe00;
			16'h9dab: y = 16'hfe00;
			16'h9dac: y = 16'hfe00;
			16'h9dad: y = 16'hfe00;
			16'h9dae: y = 16'hfe00;
			16'h9daf: y = 16'hfe00;
			16'h9db0: y = 16'hfe00;
			16'h9db1: y = 16'hfe00;
			16'h9db2: y = 16'hfe00;
			16'h9db3: y = 16'hfe00;
			16'h9db4: y = 16'hfe00;
			16'h9db5: y = 16'hfe00;
			16'h9db6: y = 16'hfe00;
			16'h9db7: y = 16'hfe00;
			16'h9db8: y = 16'hfe00;
			16'h9db9: y = 16'hfe00;
			16'h9dba: y = 16'hfe00;
			16'h9dbb: y = 16'hfe00;
			16'h9dbc: y = 16'hfe00;
			16'h9dbd: y = 16'hfe00;
			16'h9dbe: y = 16'hfe00;
			16'h9dbf: y = 16'hfe00;
			16'h9dc0: y = 16'hfe00;
			16'h9dc1: y = 16'hfe00;
			16'h9dc2: y = 16'hfe00;
			16'h9dc3: y = 16'hfe00;
			16'h9dc4: y = 16'hfe00;
			16'h9dc5: y = 16'hfe00;
			16'h9dc6: y = 16'hfe00;
			16'h9dc7: y = 16'hfe00;
			16'h9dc8: y = 16'hfe00;
			16'h9dc9: y = 16'hfe00;
			16'h9dca: y = 16'hfe00;
			16'h9dcb: y = 16'hfe00;
			16'h9dcc: y = 16'hfe00;
			16'h9dcd: y = 16'hfe00;
			16'h9dce: y = 16'hfe00;
			16'h9dcf: y = 16'hfe00;
			16'h9dd0: y = 16'hfe00;
			16'h9dd1: y = 16'hfe00;
			16'h9dd2: y = 16'hfe00;
			16'h9dd3: y = 16'hfe00;
			16'h9dd4: y = 16'hfe00;
			16'h9dd5: y = 16'hfe00;
			16'h9dd6: y = 16'hfe00;
			16'h9dd7: y = 16'hfe00;
			16'h9dd8: y = 16'hfe00;
			16'h9dd9: y = 16'hfe00;
			16'h9dda: y = 16'hfe00;
			16'h9ddb: y = 16'hfe00;
			16'h9ddc: y = 16'hfe00;
			16'h9ddd: y = 16'hfe00;
			16'h9dde: y = 16'hfe00;
			16'h9ddf: y = 16'hfe00;
			16'h9de0: y = 16'hfe00;
			16'h9de1: y = 16'hfe00;
			16'h9de2: y = 16'hfe00;
			16'h9de3: y = 16'hfe00;
			16'h9de4: y = 16'hfe00;
			16'h9de5: y = 16'hfe00;
			16'h9de6: y = 16'hfe00;
			16'h9de7: y = 16'hfe00;
			16'h9de8: y = 16'hfe00;
			16'h9de9: y = 16'hfe00;
			16'h9dea: y = 16'hfe00;
			16'h9deb: y = 16'hfe00;
			16'h9dec: y = 16'hfe00;
			16'h9ded: y = 16'hfe00;
			16'h9dee: y = 16'hfe00;
			16'h9def: y = 16'hfe00;
			16'h9df0: y = 16'hfe00;
			16'h9df1: y = 16'hfe00;
			16'h9df2: y = 16'hfe00;
			16'h9df3: y = 16'hfe00;
			16'h9df4: y = 16'hfe00;
			16'h9df5: y = 16'hfe00;
			16'h9df6: y = 16'hfe00;
			16'h9df7: y = 16'hfe00;
			16'h9df8: y = 16'hfe00;
			16'h9df9: y = 16'hfe00;
			16'h9dfa: y = 16'hfe00;
			16'h9dfb: y = 16'hfe00;
			16'h9dfc: y = 16'hfe00;
			16'h9dfd: y = 16'hfe00;
			16'h9dfe: y = 16'hfe00;
			16'h9dff: y = 16'hfe00;
			16'h9e00: y = 16'hfe00;
			16'h9e01: y = 16'hfe00;
			16'h9e02: y = 16'hfe00;
			16'h9e03: y = 16'hfe00;
			16'h9e04: y = 16'hfe00;
			16'h9e05: y = 16'hfe00;
			16'h9e06: y = 16'hfe00;
			16'h9e07: y = 16'hfe00;
			16'h9e08: y = 16'hfe00;
			16'h9e09: y = 16'hfe00;
			16'h9e0a: y = 16'hfe00;
			16'h9e0b: y = 16'hfe00;
			16'h9e0c: y = 16'hfe00;
			16'h9e0d: y = 16'hfe00;
			16'h9e0e: y = 16'hfe00;
			16'h9e0f: y = 16'hfe00;
			16'h9e10: y = 16'hfe00;
			16'h9e11: y = 16'hfe00;
			16'h9e12: y = 16'hfe00;
			16'h9e13: y = 16'hfe00;
			16'h9e14: y = 16'hfe00;
			16'h9e15: y = 16'hfe00;
			16'h9e16: y = 16'hfe00;
			16'h9e17: y = 16'hfe00;
			16'h9e18: y = 16'hfe00;
			16'h9e19: y = 16'hfe00;
			16'h9e1a: y = 16'hfe00;
			16'h9e1b: y = 16'hfe00;
			16'h9e1c: y = 16'hfe00;
			16'h9e1d: y = 16'hfe00;
			16'h9e1e: y = 16'hfe00;
			16'h9e1f: y = 16'hfe00;
			16'h9e20: y = 16'hfe00;
			16'h9e21: y = 16'hfe00;
			16'h9e22: y = 16'hfe00;
			16'h9e23: y = 16'hfe00;
			16'h9e24: y = 16'hfe00;
			16'h9e25: y = 16'hfe00;
			16'h9e26: y = 16'hfe00;
			16'h9e27: y = 16'hfe00;
			16'h9e28: y = 16'hfe00;
			16'h9e29: y = 16'hfe00;
			16'h9e2a: y = 16'hfe00;
			16'h9e2b: y = 16'hfe00;
			16'h9e2c: y = 16'hfe00;
			16'h9e2d: y = 16'hfe00;
			16'h9e2e: y = 16'hfe00;
			16'h9e2f: y = 16'hfe00;
			16'h9e30: y = 16'hfe00;
			16'h9e31: y = 16'hfe00;
			16'h9e32: y = 16'hfe00;
			16'h9e33: y = 16'hfe00;
			16'h9e34: y = 16'hfe00;
			16'h9e35: y = 16'hfe00;
			16'h9e36: y = 16'hfe00;
			16'h9e37: y = 16'hfe00;
			16'h9e38: y = 16'hfe00;
			16'h9e39: y = 16'hfe00;
			16'h9e3a: y = 16'hfe00;
			16'h9e3b: y = 16'hfe00;
			16'h9e3c: y = 16'hfe00;
			16'h9e3d: y = 16'hfe00;
			16'h9e3e: y = 16'hfe00;
			16'h9e3f: y = 16'hfe00;
			16'h9e40: y = 16'hfe00;
			16'h9e41: y = 16'hfe00;
			16'h9e42: y = 16'hfe00;
			16'h9e43: y = 16'hfe00;
			16'h9e44: y = 16'hfe00;
			16'h9e45: y = 16'hfe00;
			16'h9e46: y = 16'hfe00;
			16'h9e47: y = 16'hfe00;
			16'h9e48: y = 16'hfe00;
			16'h9e49: y = 16'hfe00;
			16'h9e4a: y = 16'hfe00;
			16'h9e4b: y = 16'hfe00;
			16'h9e4c: y = 16'hfe00;
			16'h9e4d: y = 16'hfe00;
			16'h9e4e: y = 16'hfe00;
			16'h9e4f: y = 16'hfe00;
			16'h9e50: y = 16'hfe00;
			16'h9e51: y = 16'hfe00;
			16'h9e52: y = 16'hfe00;
			16'h9e53: y = 16'hfe00;
			16'h9e54: y = 16'hfe00;
			16'h9e55: y = 16'hfe00;
			16'h9e56: y = 16'hfe00;
			16'h9e57: y = 16'hfe00;
			16'h9e58: y = 16'hfe00;
			16'h9e59: y = 16'hfe00;
			16'h9e5a: y = 16'hfe00;
			16'h9e5b: y = 16'hfe00;
			16'h9e5c: y = 16'hfe00;
			16'h9e5d: y = 16'hfe00;
			16'h9e5e: y = 16'hfe00;
			16'h9e5f: y = 16'hfe00;
			16'h9e60: y = 16'hfe00;
			16'h9e61: y = 16'hfe00;
			16'h9e62: y = 16'hfe00;
			16'h9e63: y = 16'hfe00;
			16'h9e64: y = 16'hfe00;
			16'h9e65: y = 16'hfe00;
			16'h9e66: y = 16'hfe00;
			16'h9e67: y = 16'hfe00;
			16'h9e68: y = 16'hfe00;
			16'h9e69: y = 16'hfe00;
			16'h9e6a: y = 16'hfe00;
			16'h9e6b: y = 16'hfe00;
			16'h9e6c: y = 16'hfe00;
			16'h9e6d: y = 16'hfe00;
			16'h9e6e: y = 16'hfe00;
			16'h9e6f: y = 16'hfe00;
			16'h9e70: y = 16'hfe00;
			16'h9e71: y = 16'hfe00;
			16'h9e72: y = 16'hfe00;
			16'h9e73: y = 16'hfe00;
			16'h9e74: y = 16'hfe00;
			16'h9e75: y = 16'hfe00;
			16'h9e76: y = 16'hfe00;
			16'h9e77: y = 16'hfe00;
			16'h9e78: y = 16'hfe00;
			16'h9e79: y = 16'hfe00;
			16'h9e7a: y = 16'hfe00;
			16'h9e7b: y = 16'hfe00;
			16'h9e7c: y = 16'hfe00;
			16'h9e7d: y = 16'hfe00;
			16'h9e7e: y = 16'hfe00;
			16'h9e7f: y = 16'hfe00;
			16'h9e80: y = 16'hfe00;
			16'h9e81: y = 16'hfe00;
			16'h9e82: y = 16'hfe00;
			16'h9e83: y = 16'hfe00;
			16'h9e84: y = 16'hfe00;
			16'h9e85: y = 16'hfe00;
			16'h9e86: y = 16'hfe00;
			16'h9e87: y = 16'hfe00;
			16'h9e88: y = 16'hfe00;
			16'h9e89: y = 16'hfe00;
			16'h9e8a: y = 16'hfe00;
			16'h9e8b: y = 16'hfe00;
			16'h9e8c: y = 16'hfe00;
			16'h9e8d: y = 16'hfe00;
			16'h9e8e: y = 16'hfe00;
			16'h9e8f: y = 16'hfe00;
			16'h9e90: y = 16'hfe00;
			16'h9e91: y = 16'hfe00;
			16'h9e92: y = 16'hfe00;
			16'h9e93: y = 16'hfe00;
			16'h9e94: y = 16'hfe00;
			16'h9e95: y = 16'hfe00;
			16'h9e96: y = 16'hfe00;
			16'h9e97: y = 16'hfe00;
			16'h9e98: y = 16'hfe00;
			16'h9e99: y = 16'hfe00;
			16'h9e9a: y = 16'hfe00;
			16'h9e9b: y = 16'hfe00;
			16'h9e9c: y = 16'hfe00;
			16'h9e9d: y = 16'hfe00;
			16'h9e9e: y = 16'hfe00;
			16'h9e9f: y = 16'hfe00;
			16'h9ea0: y = 16'hfe00;
			16'h9ea1: y = 16'hfe00;
			16'h9ea2: y = 16'hfe00;
			16'h9ea3: y = 16'hfe00;
			16'h9ea4: y = 16'hfe00;
			16'h9ea5: y = 16'hfe00;
			16'h9ea6: y = 16'hfe00;
			16'h9ea7: y = 16'hfe00;
			16'h9ea8: y = 16'hfe00;
			16'h9ea9: y = 16'hfe00;
			16'h9eaa: y = 16'hfe00;
			16'h9eab: y = 16'hfe00;
			16'h9eac: y = 16'hfe00;
			16'h9ead: y = 16'hfe00;
			16'h9eae: y = 16'hfe00;
			16'h9eaf: y = 16'hfe00;
			16'h9eb0: y = 16'hfe00;
			16'h9eb1: y = 16'hfe00;
			16'h9eb2: y = 16'hfe00;
			16'h9eb3: y = 16'hfe00;
			16'h9eb4: y = 16'hfe00;
			16'h9eb5: y = 16'hfe00;
			16'h9eb6: y = 16'hfe00;
			16'h9eb7: y = 16'hfe00;
			16'h9eb8: y = 16'hfe00;
			16'h9eb9: y = 16'hfe00;
			16'h9eba: y = 16'hfe00;
			16'h9ebb: y = 16'hfe00;
			16'h9ebc: y = 16'hfe00;
			16'h9ebd: y = 16'hfe00;
			16'h9ebe: y = 16'hfe00;
			16'h9ebf: y = 16'hfe00;
			16'h9ec0: y = 16'hfe00;
			16'h9ec1: y = 16'hfe00;
			16'h9ec2: y = 16'hfe00;
			16'h9ec3: y = 16'hfe00;
			16'h9ec4: y = 16'hfe00;
			16'h9ec5: y = 16'hfe00;
			16'h9ec6: y = 16'hfe00;
			16'h9ec7: y = 16'hfe00;
			16'h9ec8: y = 16'hfe00;
			16'h9ec9: y = 16'hfe00;
			16'h9eca: y = 16'hfe00;
			16'h9ecb: y = 16'hfe00;
			16'h9ecc: y = 16'hfe00;
			16'h9ecd: y = 16'hfe00;
			16'h9ece: y = 16'hfe00;
			16'h9ecf: y = 16'hfe00;
			16'h9ed0: y = 16'hfe00;
			16'h9ed1: y = 16'hfe00;
			16'h9ed2: y = 16'hfe00;
			16'h9ed3: y = 16'hfe00;
			16'h9ed4: y = 16'hfe00;
			16'h9ed5: y = 16'hfe00;
			16'h9ed6: y = 16'hfe00;
			16'h9ed7: y = 16'hfe00;
			16'h9ed8: y = 16'hfe00;
			16'h9ed9: y = 16'hfe00;
			16'h9eda: y = 16'hfe00;
			16'h9edb: y = 16'hfe00;
			16'h9edc: y = 16'hfe00;
			16'h9edd: y = 16'hfe00;
			16'h9ede: y = 16'hfe00;
			16'h9edf: y = 16'hfe00;
			16'h9ee0: y = 16'hfe00;
			16'h9ee1: y = 16'hfe00;
			16'h9ee2: y = 16'hfe00;
			16'h9ee3: y = 16'hfe00;
			16'h9ee4: y = 16'hfe00;
			16'h9ee5: y = 16'hfe00;
			16'h9ee6: y = 16'hfe00;
			16'h9ee7: y = 16'hfe00;
			16'h9ee8: y = 16'hfe00;
			16'h9ee9: y = 16'hfe00;
			16'h9eea: y = 16'hfe00;
			16'h9eeb: y = 16'hfe00;
			16'h9eec: y = 16'hfe00;
			16'h9eed: y = 16'hfe00;
			16'h9eee: y = 16'hfe00;
			16'h9eef: y = 16'hfe00;
			16'h9ef0: y = 16'hfe00;
			16'h9ef1: y = 16'hfe00;
			16'h9ef2: y = 16'hfe00;
			16'h9ef3: y = 16'hfe00;
			16'h9ef4: y = 16'hfe00;
			16'h9ef5: y = 16'hfe00;
			16'h9ef6: y = 16'hfe00;
			16'h9ef7: y = 16'hfe00;
			16'h9ef8: y = 16'hfe00;
			16'h9ef9: y = 16'hfe00;
			16'h9efa: y = 16'hfe00;
			16'h9efb: y = 16'hfe00;
			16'h9efc: y = 16'hfe00;
			16'h9efd: y = 16'hfe00;
			16'h9efe: y = 16'hfe00;
			16'h9eff: y = 16'hfe00;
			16'h9f00: y = 16'hfe00;
			16'h9f01: y = 16'hfe00;
			16'h9f02: y = 16'hfe00;
			16'h9f03: y = 16'hfe00;
			16'h9f04: y = 16'hfe00;
			16'h9f05: y = 16'hfe00;
			16'h9f06: y = 16'hfe00;
			16'h9f07: y = 16'hfe00;
			16'h9f08: y = 16'hfe00;
			16'h9f09: y = 16'hfe00;
			16'h9f0a: y = 16'hfe00;
			16'h9f0b: y = 16'hfe00;
			16'h9f0c: y = 16'hfe00;
			16'h9f0d: y = 16'hfe00;
			16'h9f0e: y = 16'hfe00;
			16'h9f0f: y = 16'hfe00;
			16'h9f10: y = 16'hfe00;
			16'h9f11: y = 16'hfe00;
			16'h9f12: y = 16'hfe00;
			16'h9f13: y = 16'hfe00;
			16'h9f14: y = 16'hfe00;
			16'h9f15: y = 16'hfe00;
			16'h9f16: y = 16'hfe00;
			16'h9f17: y = 16'hfe00;
			16'h9f18: y = 16'hfe00;
			16'h9f19: y = 16'hfe00;
			16'h9f1a: y = 16'hfe00;
			16'h9f1b: y = 16'hfe00;
			16'h9f1c: y = 16'hfe00;
			16'h9f1d: y = 16'hfe00;
			16'h9f1e: y = 16'hfe00;
			16'h9f1f: y = 16'hfe00;
			16'h9f20: y = 16'hfe00;
			16'h9f21: y = 16'hfe00;
			16'h9f22: y = 16'hfe00;
			16'h9f23: y = 16'hfe00;
			16'h9f24: y = 16'hfe00;
			16'h9f25: y = 16'hfe00;
			16'h9f26: y = 16'hfe00;
			16'h9f27: y = 16'hfe00;
			16'h9f28: y = 16'hfe00;
			16'h9f29: y = 16'hfe00;
			16'h9f2a: y = 16'hfe00;
			16'h9f2b: y = 16'hfe00;
			16'h9f2c: y = 16'hfe00;
			16'h9f2d: y = 16'hfe00;
			16'h9f2e: y = 16'hfe00;
			16'h9f2f: y = 16'hfe00;
			16'h9f30: y = 16'hfe00;
			16'h9f31: y = 16'hfe00;
			16'h9f32: y = 16'hfe00;
			16'h9f33: y = 16'hfe00;
			16'h9f34: y = 16'hfe00;
			16'h9f35: y = 16'hfe00;
			16'h9f36: y = 16'hfe00;
			16'h9f37: y = 16'hfe00;
			16'h9f38: y = 16'hfe00;
			16'h9f39: y = 16'hfe00;
			16'h9f3a: y = 16'hfe00;
			16'h9f3b: y = 16'hfe00;
			16'h9f3c: y = 16'hfe00;
			16'h9f3d: y = 16'hfe00;
			16'h9f3e: y = 16'hfe00;
			16'h9f3f: y = 16'hfe00;
			16'h9f40: y = 16'hfe00;
			16'h9f41: y = 16'hfe00;
			16'h9f42: y = 16'hfe00;
			16'h9f43: y = 16'hfe00;
			16'h9f44: y = 16'hfe00;
			16'h9f45: y = 16'hfe00;
			16'h9f46: y = 16'hfe00;
			16'h9f47: y = 16'hfe00;
			16'h9f48: y = 16'hfe00;
			16'h9f49: y = 16'hfe00;
			16'h9f4a: y = 16'hfe00;
			16'h9f4b: y = 16'hfe00;
			16'h9f4c: y = 16'hfe00;
			16'h9f4d: y = 16'hfe00;
			16'h9f4e: y = 16'hfe00;
			16'h9f4f: y = 16'hfe00;
			16'h9f50: y = 16'hfe00;
			16'h9f51: y = 16'hfe00;
			16'h9f52: y = 16'hfe00;
			16'h9f53: y = 16'hfe00;
			16'h9f54: y = 16'hfe00;
			16'h9f55: y = 16'hfe00;
			16'h9f56: y = 16'hfe00;
			16'h9f57: y = 16'hfe00;
			16'h9f58: y = 16'hfe00;
			16'h9f59: y = 16'hfe00;
			16'h9f5a: y = 16'hfe00;
			16'h9f5b: y = 16'hfe00;
			16'h9f5c: y = 16'hfe00;
			16'h9f5d: y = 16'hfe00;
			16'h9f5e: y = 16'hfe00;
			16'h9f5f: y = 16'hfe00;
			16'h9f60: y = 16'hfe00;
			16'h9f61: y = 16'hfe00;
			16'h9f62: y = 16'hfe00;
			16'h9f63: y = 16'hfe00;
			16'h9f64: y = 16'hfe00;
			16'h9f65: y = 16'hfe00;
			16'h9f66: y = 16'hfe00;
			16'h9f67: y = 16'hfe00;
			16'h9f68: y = 16'hfe00;
			16'h9f69: y = 16'hfe00;
			16'h9f6a: y = 16'hfe00;
			16'h9f6b: y = 16'hfe00;
			16'h9f6c: y = 16'hfe00;
			16'h9f6d: y = 16'hfe00;
			16'h9f6e: y = 16'hfe00;
			16'h9f6f: y = 16'hfe00;
			16'h9f70: y = 16'hfe00;
			16'h9f71: y = 16'hfe00;
			16'h9f72: y = 16'hfe00;
			16'h9f73: y = 16'hfe00;
			16'h9f74: y = 16'hfe00;
			16'h9f75: y = 16'hfe00;
			16'h9f76: y = 16'hfe00;
			16'h9f77: y = 16'hfe00;
			16'h9f78: y = 16'hfe00;
			16'h9f79: y = 16'hfe00;
			16'h9f7a: y = 16'hfe00;
			16'h9f7b: y = 16'hfe00;
			16'h9f7c: y = 16'hfe00;
			16'h9f7d: y = 16'hfe00;
			16'h9f7e: y = 16'hfe00;
			16'h9f7f: y = 16'hfe00;
			16'h9f80: y = 16'hfe00;
			16'h9f81: y = 16'hfe00;
			16'h9f82: y = 16'hfe00;
			16'h9f83: y = 16'hfe00;
			16'h9f84: y = 16'hfe00;
			16'h9f85: y = 16'hfe00;
			16'h9f86: y = 16'hfe00;
			16'h9f87: y = 16'hfe00;
			16'h9f88: y = 16'hfe00;
			16'h9f89: y = 16'hfe00;
			16'h9f8a: y = 16'hfe00;
			16'h9f8b: y = 16'hfe00;
			16'h9f8c: y = 16'hfe00;
			16'h9f8d: y = 16'hfe00;
			16'h9f8e: y = 16'hfe00;
			16'h9f8f: y = 16'hfe00;
			16'h9f90: y = 16'hfe00;
			16'h9f91: y = 16'hfe00;
			16'h9f92: y = 16'hfe00;
			16'h9f93: y = 16'hfe00;
			16'h9f94: y = 16'hfe00;
			16'h9f95: y = 16'hfe00;
			16'h9f96: y = 16'hfe00;
			16'h9f97: y = 16'hfe00;
			16'h9f98: y = 16'hfe00;
			16'h9f99: y = 16'hfe00;
			16'h9f9a: y = 16'hfe00;
			16'h9f9b: y = 16'hfe00;
			16'h9f9c: y = 16'hfe00;
			16'h9f9d: y = 16'hfe00;
			16'h9f9e: y = 16'hfe00;
			16'h9f9f: y = 16'hfe00;
			16'h9fa0: y = 16'hfe00;
			16'h9fa1: y = 16'hfe00;
			16'h9fa2: y = 16'hfe00;
			16'h9fa3: y = 16'hfe00;
			16'h9fa4: y = 16'hfe00;
			16'h9fa5: y = 16'hfe00;
			16'h9fa6: y = 16'hfe00;
			16'h9fa7: y = 16'hfe00;
			16'h9fa8: y = 16'hfe00;
			16'h9fa9: y = 16'hfe00;
			16'h9faa: y = 16'hfe00;
			16'h9fab: y = 16'hfe00;
			16'h9fac: y = 16'hfe00;
			16'h9fad: y = 16'hfe00;
			16'h9fae: y = 16'hfe00;
			16'h9faf: y = 16'hfe00;
			16'h9fb0: y = 16'hfe00;
			16'h9fb1: y = 16'hfe00;
			16'h9fb2: y = 16'hfe00;
			16'h9fb3: y = 16'hfe00;
			16'h9fb4: y = 16'hfe00;
			16'h9fb5: y = 16'hfe00;
			16'h9fb6: y = 16'hfe00;
			16'h9fb7: y = 16'hfe00;
			16'h9fb8: y = 16'hfe00;
			16'h9fb9: y = 16'hfe00;
			16'h9fba: y = 16'hfe00;
			16'h9fbb: y = 16'hfe00;
			16'h9fbc: y = 16'hfe00;
			16'h9fbd: y = 16'hfe00;
			16'h9fbe: y = 16'hfe00;
			16'h9fbf: y = 16'hfe00;
			16'h9fc0: y = 16'hfe00;
			16'h9fc1: y = 16'hfe00;
			16'h9fc2: y = 16'hfe00;
			16'h9fc3: y = 16'hfe00;
			16'h9fc4: y = 16'hfe00;
			16'h9fc5: y = 16'hfe00;
			16'h9fc6: y = 16'hfe00;
			16'h9fc7: y = 16'hfe00;
			16'h9fc8: y = 16'hfe00;
			16'h9fc9: y = 16'hfe00;
			16'h9fca: y = 16'hfe00;
			16'h9fcb: y = 16'hfe00;
			16'h9fcc: y = 16'hfe00;
			16'h9fcd: y = 16'hfe00;
			16'h9fce: y = 16'hfe00;
			16'h9fcf: y = 16'hfe00;
			16'h9fd0: y = 16'hfe00;
			16'h9fd1: y = 16'hfe00;
			16'h9fd2: y = 16'hfe00;
			16'h9fd3: y = 16'hfe00;
			16'h9fd4: y = 16'hfe00;
			16'h9fd5: y = 16'hfe00;
			16'h9fd6: y = 16'hfe00;
			16'h9fd7: y = 16'hfe00;
			16'h9fd8: y = 16'hfe00;
			16'h9fd9: y = 16'hfe00;
			16'h9fda: y = 16'hfe00;
			16'h9fdb: y = 16'hfe00;
			16'h9fdc: y = 16'hfe00;
			16'h9fdd: y = 16'hfe00;
			16'h9fde: y = 16'hfe00;
			16'h9fdf: y = 16'hfe00;
			16'h9fe0: y = 16'hfe00;
			16'h9fe1: y = 16'hfe00;
			16'h9fe2: y = 16'hfe00;
			16'h9fe3: y = 16'hfe00;
			16'h9fe4: y = 16'hfe00;
			16'h9fe5: y = 16'hfe00;
			16'h9fe6: y = 16'hfe00;
			16'h9fe7: y = 16'hfe00;
			16'h9fe8: y = 16'hfe00;
			16'h9fe9: y = 16'hfe00;
			16'h9fea: y = 16'hfe00;
			16'h9feb: y = 16'hfe00;
			16'h9fec: y = 16'hfe00;
			16'h9fed: y = 16'hfe00;
			16'h9fee: y = 16'hfe00;
			16'h9fef: y = 16'hfe00;
			16'h9ff0: y = 16'hfe00;
			16'h9ff1: y = 16'hfe00;
			16'h9ff2: y = 16'hfe00;
			16'h9ff3: y = 16'hfe00;
			16'h9ff4: y = 16'hfe00;
			16'h9ff5: y = 16'hfe00;
			16'h9ff6: y = 16'hfe00;
			16'h9ff7: y = 16'hfe00;
			16'h9ff8: y = 16'hfe00;
			16'h9ff9: y = 16'hfe00;
			16'h9ffa: y = 16'hfe00;
			16'h9ffb: y = 16'hfe00;
			16'h9ffc: y = 16'hfe00;
			16'h9ffd: y = 16'hfe00;
			16'h9ffe: y = 16'hfe00;
			16'h9fff: y = 16'hfe00;
			16'ha000: y = 16'hfe00;
			16'ha001: y = 16'hfe00;
			16'ha002: y = 16'hfe00;
			16'ha003: y = 16'hfe00;
			16'ha004: y = 16'hfe00;
			16'ha005: y = 16'hfe00;
			16'ha006: y = 16'hfe00;
			16'ha007: y = 16'hfe00;
			16'ha008: y = 16'hfe00;
			16'ha009: y = 16'hfe00;
			16'ha00a: y = 16'hfe00;
			16'ha00b: y = 16'hfe00;
			16'ha00c: y = 16'hfe00;
			16'ha00d: y = 16'hfe00;
			16'ha00e: y = 16'hfe00;
			16'ha00f: y = 16'hfe00;
			16'ha010: y = 16'hfe00;
			16'ha011: y = 16'hfe00;
			16'ha012: y = 16'hfe00;
			16'ha013: y = 16'hfe00;
			16'ha014: y = 16'hfe00;
			16'ha015: y = 16'hfe00;
			16'ha016: y = 16'hfe00;
			16'ha017: y = 16'hfe00;
			16'ha018: y = 16'hfe00;
			16'ha019: y = 16'hfe00;
			16'ha01a: y = 16'hfe00;
			16'ha01b: y = 16'hfe00;
			16'ha01c: y = 16'hfe00;
			16'ha01d: y = 16'hfe00;
			16'ha01e: y = 16'hfe00;
			16'ha01f: y = 16'hfe00;
			16'ha020: y = 16'hfe00;
			16'ha021: y = 16'hfe00;
			16'ha022: y = 16'hfe00;
			16'ha023: y = 16'hfe00;
			16'ha024: y = 16'hfe00;
			16'ha025: y = 16'hfe00;
			16'ha026: y = 16'hfe00;
			16'ha027: y = 16'hfe00;
			16'ha028: y = 16'hfe00;
			16'ha029: y = 16'hfe00;
			16'ha02a: y = 16'hfe00;
			16'ha02b: y = 16'hfe00;
			16'ha02c: y = 16'hfe00;
			16'ha02d: y = 16'hfe00;
			16'ha02e: y = 16'hfe00;
			16'ha02f: y = 16'hfe00;
			16'ha030: y = 16'hfe00;
			16'ha031: y = 16'hfe00;
			16'ha032: y = 16'hfe00;
			16'ha033: y = 16'hfe00;
			16'ha034: y = 16'hfe00;
			16'ha035: y = 16'hfe00;
			16'ha036: y = 16'hfe00;
			16'ha037: y = 16'hfe00;
			16'ha038: y = 16'hfe00;
			16'ha039: y = 16'hfe00;
			16'ha03a: y = 16'hfe00;
			16'ha03b: y = 16'hfe00;
			16'ha03c: y = 16'hfe00;
			16'ha03d: y = 16'hfe00;
			16'ha03e: y = 16'hfe00;
			16'ha03f: y = 16'hfe00;
			16'ha040: y = 16'hfe00;
			16'ha041: y = 16'hfe00;
			16'ha042: y = 16'hfe00;
			16'ha043: y = 16'hfe00;
			16'ha044: y = 16'hfe00;
			16'ha045: y = 16'hfe00;
			16'ha046: y = 16'hfe00;
			16'ha047: y = 16'hfe00;
			16'ha048: y = 16'hfe00;
			16'ha049: y = 16'hfe00;
			16'ha04a: y = 16'hfe00;
			16'ha04b: y = 16'hfe00;
			16'ha04c: y = 16'hfe00;
			16'ha04d: y = 16'hfe00;
			16'ha04e: y = 16'hfe00;
			16'ha04f: y = 16'hfe00;
			16'ha050: y = 16'hfe00;
			16'ha051: y = 16'hfe00;
			16'ha052: y = 16'hfe00;
			16'ha053: y = 16'hfe00;
			16'ha054: y = 16'hfe00;
			16'ha055: y = 16'hfe00;
			16'ha056: y = 16'hfe00;
			16'ha057: y = 16'hfe00;
			16'ha058: y = 16'hfe00;
			16'ha059: y = 16'hfe00;
			16'ha05a: y = 16'hfe00;
			16'ha05b: y = 16'hfe00;
			16'ha05c: y = 16'hfe00;
			16'ha05d: y = 16'hfe00;
			16'ha05e: y = 16'hfe00;
			16'ha05f: y = 16'hfe00;
			16'ha060: y = 16'hfe00;
			16'ha061: y = 16'hfe00;
			16'ha062: y = 16'hfe00;
			16'ha063: y = 16'hfe00;
			16'ha064: y = 16'hfe00;
			16'ha065: y = 16'hfe00;
			16'ha066: y = 16'hfe00;
			16'ha067: y = 16'hfe00;
			16'ha068: y = 16'hfe00;
			16'ha069: y = 16'hfe00;
			16'ha06a: y = 16'hfe00;
			16'ha06b: y = 16'hfe00;
			16'ha06c: y = 16'hfe00;
			16'ha06d: y = 16'hfe00;
			16'ha06e: y = 16'hfe00;
			16'ha06f: y = 16'hfe00;
			16'ha070: y = 16'hfe00;
			16'ha071: y = 16'hfe00;
			16'ha072: y = 16'hfe00;
			16'ha073: y = 16'hfe00;
			16'ha074: y = 16'hfe00;
			16'ha075: y = 16'hfe00;
			16'ha076: y = 16'hfe00;
			16'ha077: y = 16'hfe00;
			16'ha078: y = 16'hfe00;
			16'ha079: y = 16'hfe00;
			16'ha07a: y = 16'hfe00;
			16'ha07b: y = 16'hfe00;
			16'ha07c: y = 16'hfe00;
			16'ha07d: y = 16'hfe00;
			16'ha07e: y = 16'hfe00;
			16'ha07f: y = 16'hfe00;
			16'ha080: y = 16'hfe00;
			16'ha081: y = 16'hfe00;
			16'ha082: y = 16'hfe00;
			16'ha083: y = 16'hfe00;
			16'ha084: y = 16'hfe00;
			16'ha085: y = 16'hfe00;
			16'ha086: y = 16'hfe00;
			16'ha087: y = 16'hfe00;
			16'ha088: y = 16'hfe00;
			16'ha089: y = 16'hfe00;
			16'ha08a: y = 16'hfe00;
			16'ha08b: y = 16'hfe00;
			16'ha08c: y = 16'hfe00;
			16'ha08d: y = 16'hfe00;
			16'ha08e: y = 16'hfe00;
			16'ha08f: y = 16'hfe00;
			16'ha090: y = 16'hfe00;
			16'ha091: y = 16'hfe00;
			16'ha092: y = 16'hfe00;
			16'ha093: y = 16'hfe00;
			16'ha094: y = 16'hfe00;
			16'ha095: y = 16'hfe00;
			16'ha096: y = 16'hfe00;
			16'ha097: y = 16'hfe00;
			16'ha098: y = 16'hfe00;
			16'ha099: y = 16'hfe00;
			16'ha09a: y = 16'hfe00;
			16'ha09b: y = 16'hfe00;
			16'ha09c: y = 16'hfe00;
			16'ha09d: y = 16'hfe00;
			16'ha09e: y = 16'hfe00;
			16'ha09f: y = 16'hfe00;
			16'ha0a0: y = 16'hfe00;
			16'ha0a1: y = 16'hfe00;
			16'ha0a2: y = 16'hfe00;
			16'ha0a3: y = 16'hfe00;
			16'ha0a4: y = 16'hfe00;
			16'ha0a5: y = 16'hfe00;
			16'ha0a6: y = 16'hfe00;
			16'ha0a7: y = 16'hfe00;
			16'ha0a8: y = 16'hfe00;
			16'ha0a9: y = 16'hfe00;
			16'ha0aa: y = 16'hfe00;
			16'ha0ab: y = 16'hfe00;
			16'ha0ac: y = 16'hfe00;
			16'ha0ad: y = 16'hfe00;
			16'ha0ae: y = 16'hfe00;
			16'ha0af: y = 16'hfe00;
			16'ha0b0: y = 16'hfe00;
			16'ha0b1: y = 16'hfe00;
			16'ha0b2: y = 16'hfe00;
			16'ha0b3: y = 16'hfe00;
			16'ha0b4: y = 16'hfe00;
			16'ha0b5: y = 16'hfe00;
			16'ha0b6: y = 16'hfe00;
			16'ha0b7: y = 16'hfe00;
			16'ha0b8: y = 16'hfe00;
			16'ha0b9: y = 16'hfe00;
			16'ha0ba: y = 16'hfe00;
			16'ha0bb: y = 16'hfe00;
			16'ha0bc: y = 16'hfe00;
			16'ha0bd: y = 16'hfe00;
			16'ha0be: y = 16'hfe00;
			16'ha0bf: y = 16'hfe00;
			16'ha0c0: y = 16'hfe00;
			16'ha0c1: y = 16'hfe00;
			16'ha0c2: y = 16'hfe00;
			16'ha0c3: y = 16'hfe00;
			16'ha0c4: y = 16'hfe00;
			16'ha0c5: y = 16'hfe00;
			16'ha0c6: y = 16'hfe00;
			16'ha0c7: y = 16'hfe00;
			16'ha0c8: y = 16'hfe00;
			16'ha0c9: y = 16'hfe00;
			16'ha0ca: y = 16'hfe00;
			16'ha0cb: y = 16'hfe00;
			16'ha0cc: y = 16'hfe00;
			16'ha0cd: y = 16'hfe00;
			16'ha0ce: y = 16'hfe00;
			16'ha0cf: y = 16'hfe00;
			16'ha0d0: y = 16'hfe00;
			16'ha0d1: y = 16'hfe00;
			16'ha0d2: y = 16'hfe00;
			16'ha0d3: y = 16'hfe00;
			16'ha0d4: y = 16'hfe00;
			16'ha0d5: y = 16'hfe00;
			16'ha0d6: y = 16'hfe00;
			16'ha0d7: y = 16'hfe00;
			16'ha0d8: y = 16'hfe00;
			16'ha0d9: y = 16'hfe00;
			16'ha0da: y = 16'hfe00;
			16'ha0db: y = 16'hfe00;
			16'ha0dc: y = 16'hfe00;
			16'ha0dd: y = 16'hfe00;
			16'ha0de: y = 16'hfe00;
			16'ha0df: y = 16'hfe00;
			16'ha0e0: y = 16'hfe00;
			16'ha0e1: y = 16'hfe00;
			16'ha0e2: y = 16'hfe00;
			16'ha0e3: y = 16'hfe00;
			16'ha0e4: y = 16'hfe00;
			16'ha0e5: y = 16'hfe00;
			16'ha0e6: y = 16'hfe00;
			16'ha0e7: y = 16'hfe00;
			16'ha0e8: y = 16'hfe00;
			16'ha0e9: y = 16'hfe00;
			16'ha0ea: y = 16'hfe00;
			16'ha0eb: y = 16'hfe00;
			16'ha0ec: y = 16'hfe00;
			16'ha0ed: y = 16'hfe00;
			16'ha0ee: y = 16'hfe00;
			16'ha0ef: y = 16'hfe00;
			16'ha0f0: y = 16'hfe00;
			16'ha0f1: y = 16'hfe00;
			16'ha0f2: y = 16'hfe00;
			16'ha0f3: y = 16'hfe00;
			16'ha0f4: y = 16'hfe00;
			16'ha0f5: y = 16'hfe00;
			16'ha0f6: y = 16'hfe00;
			16'ha0f7: y = 16'hfe00;
			16'ha0f8: y = 16'hfe00;
			16'ha0f9: y = 16'hfe00;
			16'ha0fa: y = 16'hfe00;
			16'ha0fb: y = 16'hfe00;
			16'ha0fc: y = 16'hfe00;
			16'ha0fd: y = 16'hfe00;
			16'ha0fe: y = 16'hfe00;
			16'ha0ff: y = 16'hfe00;
			16'ha100: y = 16'hfe00;
			16'ha101: y = 16'hfe00;
			16'ha102: y = 16'hfe00;
			16'ha103: y = 16'hfe00;
			16'ha104: y = 16'hfe00;
			16'ha105: y = 16'hfe00;
			16'ha106: y = 16'hfe00;
			16'ha107: y = 16'hfe00;
			16'ha108: y = 16'hfe00;
			16'ha109: y = 16'hfe00;
			16'ha10a: y = 16'hfe00;
			16'ha10b: y = 16'hfe00;
			16'ha10c: y = 16'hfe00;
			16'ha10d: y = 16'hfe00;
			16'ha10e: y = 16'hfe00;
			16'ha10f: y = 16'hfe00;
			16'ha110: y = 16'hfe00;
			16'ha111: y = 16'hfe00;
			16'ha112: y = 16'hfe00;
			16'ha113: y = 16'hfe00;
			16'ha114: y = 16'hfe00;
			16'ha115: y = 16'hfe00;
			16'ha116: y = 16'hfe00;
			16'ha117: y = 16'hfe00;
			16'ha118: y = 16'hfe00;
			16'ha119: y = 16'hfe00;
			16'ha11a: y = 16'hfe00;
			16'ha11b: y = 16'hfe00;
			16'ha11c: y = 16'hfe00;
			16'ha11d: y = 16'hfe00;
			16'ha11e: y = 16'hfe00;
			16'ha11f: y = 16'hfe00;
			16'ha120: y = 16'hfe00;
			16'ha121: y = 16'hfe00;
			16'ha122: y = 16'hfe00;
			16'ha123: y = 16'hfe00;
			16'ha124: y = 16'hfe00;
			16'ha125: y = 16'hfe00;
			16'ha126: y = 16'hfe00;
			16'ha127: y = 16'hfe00;
			16'ha128: y = 16'hfe00;
			16'ha129: y = 16'hfe00;
			16'ha12a: y = 16'hfe00;
			16'ha12b: y = 16'hfe00;
			16'ha12c: y = 16'hfe00;
			16'ha12d: y = 16'hfe00;
			16'ha12e: y = 16'hfe00;
			16'ha12f: y = 16'hfe00;
			16'ha130: y = 16'hfe00;
			16'ha131: y = 16'hfe00;
			16'ha132: y = 16'hfe00;
			16'ha133: y = 16'hfe00;
			16'ha134: y = 16'hfe00;
			16'ha135: y = 16'hfe00;
			16'ha136: y = 16'hfe00;
			16'ha137: y = 16'hfe00;
			16'ha138: y = 16'hfe00;
			16'ha139: y = 16'hfe00;
			16'ha13a: y = 16'hfe00;
			16'ha13b: y = 16'hfe00;
			16'ha13c: y = 16'hfe00;
			16'ha13d: y = 16'hfe00;
			16'ha13e: y = 16'hfe00;
			16'ha13f: y = 16'hfe00;
			16'ha140: y = 16'hfe00;
			16'ha141: y = 16'hfe00;
			16'ha142: y = 16'hfe00;
			16'ha143: y = 16'hfe00;
			16'ha144: y = 16'hfe00;
			16'ha145: y = 16'hfe00;
			16'ha146: y = 16'hfe00;
			16'ha147: y = 16'hfe00;
			16'ha148: y = 16'hfe00;
			16'ha149: y = 16'hfe00;
			16'ha14a: y = 16'hfe00;
			16'ha14b: y = 16'hfe00;
			16'ha14c: y = 16'hfe00;
			16'ha14d: y = 16'hfe00;
			16'ha14e: y = 16'hfe00;
			16'ha14f: y = 16'hfe00;
			16'ha150: y = 16'hfe00;
			16'ha151: y = 16'hfe00;
			16'ha152: y = 16'hfe00;
			16'ha153: y = 16'hfe00;
			16'ha154: y = 16'hfe00;
			16'ha155: y = 16'hfe00;
			16'ha156: y = 16'hfe00;
			16'ha157: y = 16'hfe00;
			16'ha158: y = 16'hfe00;
			16'ha159: y = 16'hfe00;
			16'ha15a: y = 16'hfe00;
			16'ha15b: y = 16'hfe00;
			16'ha15c: y = 16'hfe00;
			16'ha15d: y = 16'hfe00;
			16'ha15e: y = 16'hfe00;
			16'ha15f: y = 16'hfe00;
			16'ha160: y = 16'hfe00;
			16'ha161: y = 16'hfe00;
			16'ha162: y = 16'hfe00;
			16'ha163: y = 16'hfe00;
			16'ha164: y = 16'hfe00;
			16'ha165: y = 16'hfe00;
			16'ha166: y = 16'hfe00;
			16'ha167: y = 16'hfe00;
			16'ha168: y = 16'hfe00;
			16'ha169: y = 16'hfe00;
			16'ha16a: y = 16'hfe00;
			16'ha16b: y = 16'hfe00;
			16'ha16c: y = 16'hfe00;
			16'ha16d: y = 16'hfe00;
			16'ha16e: y = 16'hfe00;
			16'ha16f: y = 16'hfe00;
			16'ha170: y = 16'hfe00;
			16'ha171: y = 16'hfe00;
			16'ha172: y = 16'hfe00;
			16'ha173: y = 16'hfe00;
			16'ha174: y = 16'hfe00;
			16'ha175: y = 16'hfe00;
			16'ha176: y = 16'hfe00;
			16'ha177: y = 16'hfe00;
			16'ha178: y = 16'hfe00;
			16'ha179: y = 16'hfe00;
			16'ha17a: y = 16'hfe00;
			16'ha17b: y = 16'hfe00;
			16'ha17c: y = 16'hfe00;
			16'ha17d: y = 16'hfe00;
			16'ha17e: y = 16'hfe00;
			16'ha17f: y = 16'hfe00;
			16'ha180: y = 16'hfe00;
			16'ha181: y = 16'hfe00;
			16'ha182: y = 16'hfe00;
			16'ha183: y = 16'hfe00;
			16'ha184: y = 16'hfe00;
			16'ha185: y = 16'hfe00;
			16'ha186: y = 16'hfe00;
			16'ha187: y = 16'hfe00;
			16'ha188: y = 16'hfe00;
			16'ha189: y = 16'hfe00;
			16'ha18a: y = 16'hfe00;
			16'ha18b: y = 16'hfe00;
			16'ha18c: y = 16'hfe00;
			16'ha18d: y = 16'hfe00;
			16'ha18e: y = 16'hfe00;
			16'ha18f: y = 16'hfe00;
			16'ha190: y = 16'hfe00;
			16'ha191: y = 16'hfe00;
			16'ha192: y = 16'hfe00;
			16'ha193: y = 16'hfe00;
			16'ha194: y = 16'hfe00;
			16'ha195: y = 16'hfe00;
			16'ha196: y = 16'hfe00;
			16'ha197: y = 16'hfe00;
			16'ha198: y = 16'hfe00;
			16'ha199: y = 16'hfe00;
			16'ha19a: y = 16'hfe00;
			16'ha19b: y = 16'hfe00;
			16'ha19c: y = 16'hfe00;
			16'ha19d: y = 16'hfe00;
			16'ha19e: y = 16'hfe00;
			16'ha19f: y = 16'hfe00;
			16'ha1a0: y = 16'hfe00;
			16'ha1a1: y = 16'hfe00;
			16'ha1a2: y = 16'hfe00;
			16'ha1a3: y = 16'hfe00;
			16'ha1a4: y = 16'hfe00;
			16'ha1a5: y = 16'hfe00;
			16'ha1a6: y = 16'hfe00;
			16'ha1a7: y = 16'hfe00;
			16'ha1a8: y = 16'hfe00;
			16'ha1a9: y = 16'hfe00;
			16'ha1aa: y = 16'hfe00;
			16'ha1ab: y = 16'hfe00;
			16'ha1ac: y = 16'hfe00;
			16'ha1ad: y = 16'hfe00;
			16'ha1ae: y = 16'hfe00;
			16'ha1af: y = 16'hfe00;
			16'ha1b0: y = 16'hfe00;
			16'ha1b1: y = 16'hfe00;
			16'ha1b2: y = 16'hfe00;
			16'ha1b3: y = 16'hfe00;
			16'ha1b4: y = 16'hfe00;
			16'ha1b5: y = 16'hfe00;
			16'ha1b6: y = 16'hfe00;
			16'ha1b7: y = 16'hfe00;
			16'ha1b8: y = 16'hfe00;
			16'ha1b9: y = 16'hfe00;
			16'ha1ba: y = 16'hfe00;
			16'ha1bb: y = 16'hfe00;
			16'ha1bc: y = 16'hfe00;
			16'ha1bd: y = 16'hfe00;
			16'ha1be: y = 16'hfe00;
			16'ha1bf: y = 16'hfe00;
			16'ha1c0: y = 16'hfe00;
			16'ha1c1: y = 16'hfe00;
			16'ha1c2: y = 16'hfe00;
			16'ha1c3: y = 16'hfe00;
			16'ha1c4: y = 16'hfe00;
			16'ha1c5: y = 16'hfe00;
			16'ha1c6: y = 16'hfe00;
			16'ha1c7: y = 16'hfe00;
			16'ha1c8: y = 16'hfe00;
			16'ha1c9: y = 16'hfe00;
			16'ha1ca: y = 16'hfe00;
			16'ha1cb: y = 16'hfe00;
			16'ha1cc: y = 16'hfe00;
			16'ha1cd: y = 16'hfe00;
			16'ha1ce: y = 16'hfe00;
			16'ha1cf: y = 16'hfe00;
			16'ha1d0: y = 16'hfe00;
			16'ha1d1: y = 16'hfe00;
			16'ha1d2: y = 16'hfe00;
			16'ha1d3: y = 16'hfe00;
			16'ha1d4: y = 16'hfe00;
			16'ha1d5: y = 16'hfe00;
			16'ha1d6: y = 16'hfe00;
			16'ha1d7: y = 16'hfe00;
			16'ha1d8: y = 16'hfe00;
			16'ha1d9: y = 16'hfe00;
			16'ha1da: y = 16'hfe00;
			16'ha1db: y = 16'hfe00;
			16'ha1dc: y = 16'hfe00;
			16'ha1dd: y = 16'hfe00;
			16'ha1de: y = 16'hfe00;
			16'ha1df: y = 16'hfe00;
			16'ha1e0: y = 16'hfe00;
			16'ha1e1: y = 16'hfe00;
			16'ha1e2: y = 16'hfe00;
			16'ha1e3: y = 16'hfe00;
			16'ha1e4: y = 16'hfe00;
			16'ha1e5: y = 16'hfe00;
			16'ha1e6: y = 16'hfe00;
			16'ha1e7: y = 16'hfe00;
			16'ha1e8: y = 16'hfe00;
			16'ha1e9: y = 16'hfe00;
			16'ha1ea: y = 16'hfe00;
			16'ha1eb: y = 16'hfe00;
			16'ha1ec: y = 16'hfe00;
			16'ha1ed: y = 16'hfe00;
			16'ha1ee: y = 16'hfe00;
			16'ha1ef: y = 16'hfe00;
			16'ha1f0: y = 16'hfe00;
			16'ha1f1: y = 16'hfe00;
			16'ha1f2: y = 16'hfe00;
			16'ha1f3: y = 16'hfe00;
			16'ha1f4: y = 16'hfe00;
			16'ha1f5: y = 16'hfe00;
			16'ha1f6: y = 16'hfe00;
			16'ha1f7: y = 16'hfe00;
			16'ha1f8: y = 16'hfe00;
			16'ha1f9: y = 16'hfe00;
			16'ha1fa: y = 16'hfe00;
			16'ha1fb: y = 16'hfe00;
			16'ha1fc: y = 16'hfe00;
			16'ha1fd: y = 16'hfe00;
			16'ha1fe: y = 16'hfe00;
			16'ha1ff: y = 16'hfe00;
			16'ha200: y = 16'hfe00;
			16'ha201: y = 16'hfe00;
			16'ha202: y = 16'hfe00;
			16'ha203: y = 16'hfe00;
			16'ha204: y = 16'hfe00;
			16'ha205: y = 16'hfe00;
			16'ha206: y = 16'hfe00;
			16'ha207: y = 16'hfe00;
			16'ha208: y = 16'hfe00;
			16'ha209: y = 16'hfe00;
			16'ha20a: y = 16'hfe00;
			16'ha20b: y = 16'hfe00;
			16'ha20c: y = 16'hfe00;
			16'ha20d: y = 16'hfe00;
			16'ha20e: y = 16'hfe00;
			16'ha20f: y = 16'hfe00;
			16'ha210: y = 16'hfe00;
			16'ha211: y = 16'hfe00;
			16'ha212: y = 16'hfe00;
			16'ha213: y = 16'hfe00;
			16'ha214: y = 16'hfe00;
			16'ha215: y = 16'hfe00;
			16'ha216: y = 16'hfe00;
			16'ha217: y = 16'hfe00;
			16'ha218: y = 16'hfe00;
			16'ha219: y = 16'hfe00;
			16'ha21a: y = 16'hfe00;
			16'ha21b: y = 16'hfe00;
			16'ha21c: y = 16'hfe00;
			16'ha21d: y = 16'hfe00;
			16'ha21e: y = 16'hfe00;
			16'ha21f: y = 16'hfe00;
			16'ha220: y = 16'hfe00;
			16'ha221: y = 16'hfe00;
			16'ha222: y = 16'hfe00;
			16'ha223: y = 16'hfe00;
			16'ha224: y = 16'hfe00;
			16'ha225: y = 16'hfe00;
			16'ha226: y = 16'hfe00;
			16'ha227: y = 16'hfe00;
			16'ha228: y = 16'hfe00;
			16'ha229: y = 16'hfe00;
			16'ha22a: y = 16'hfe00;
			16'ha22b: y = 16'hfe00;
			16'ha22c: y = 16'hfe00;
			16'ha22d: y = 16'hfe00;
			16'ha22e: y = 16'hfe00;
			16'ha22f: y = 16'hfe00;
			16'ha230: y = 16'hfe00;
			16'ha231: y = 16'hfe00;
			16'ha232: y = 16'hfe00;
			16'ha233: y = 16'hfe00;
			16'ha234: y = 16'hfe00;
			16'ha235: y = 16'hfe00;
			16'ha236: y = 16'hfe00;
			16'ha237: y = 16'hfe00;
			16'ha238: y = 16'hfe00;
			16'ha239: y = 16'hfe00;
			16'ha23a: y = 16'hfe00;
			16'ha23b: y = 16'hfe00;
			16'ha23c: y = 16'hfe00;
			16'ha23d: y = 16'hfe00;
			16'ha23e: y = 16'hfe00;
			16'ha23f: y = 16'hfe00;
			16'ha240: y = 16'hfe00;
			16'ha241: y = 16'hfe00;
			16'ha242: y = 16'hfe00;
			16'ha243: y = 16'hfe00;
			16'ha244: y = 16'hfe00;
			16'ha245: y = 16'hfe00;
			16'ha246: y = 16'hfe00;
			16'ha247: y = 16'hfe00;
			16'ha248: y = 16'hfe00;
			16'ha249: y = 16'hfe00;
			16'ha24a: y = 16'hfe00;
			16'ha24b: y = 16'hfe00;
			16'ha24c: y = 16'hfe00;
			16'ha24d: y = 16'hfe00;
			16'ha24e: y = 16'hfe00;
			16'ha24f: y = 16'hfe00;
			16'ha250: y = 16'hfe00;
			16'ha251: y = 16'hfe00;
			16'ha252: y = 16'hfe00;
			16'ha253: y = 16'hfe00;
			16'ha254: y = 16'hfe00;
			16'ha255: y = 16'hfe00;
			16'ha256: y = 16'hfe00;
			16'ha257: y = 16'hfe00;
			16'ha258: y = 16'hfe00;
			16'ha259: y = 16'hfe00;
			16'ha25a: y = 16'hfe00;
			16'ha25b: y = 16'hfe00;
			16'ha25c: y = 16'hfe00;
			16'ha25d: y = 16'hfe00;
			16'ha25e: y = 16'hfe00;
			16'ha25f: y = 16'hfe00;
			16'ha260: y = 16'hfe00;
			16'ha261: y = 16'hfe00;
			16'ha262: y = 16'hfe00;
			16'ha263: y = 16'hfe00;
			16'ha264: y = 16'hfe00;
			16'ha265: y = 16'hfe00;
			16'ha266: y = 16'hfe00;
			16'ha267: y = 16'hfe00;
			16'ha268: y = 16'hfe00;
			16'ha269: y = 16'hfe00;
			16'ha26a: y = 16'hfe00;
			16'ha26b: y = 16'hfe00;
			16'ha26c: y = 16'hfe00;
			16'ha26d: y = 16'hfe00;
			16'ha26e: y = 16'hfe00;
			16'ha26f: y = 16'hfe00;
			16'ha270: y = 16'hfe00;
			16'ha271: y = 16'hfe00;
			16'ha272: y = 16'hfe00;
			16'ha273: y = 16'hfe00;
			16'ha274: y = 16'hfe00;
			16'ha275: y = 16'hfe00;
			16'ha276: y = 16'hfe00;
			16'ha277: y = 16'hfe00;
			16'ha278: y = 16'hfe00;
			16'ha279: y = 16'hfe00;
			16'ha27a: y = 16'hfe00;
			16'ha27b: y = 16'hfe00;
			16'ha27c: y = 16'hfe00;
			16'ha27d: y = 16'hfe00;
			16'ha27e: y = 16'hfe00;
			16'ha27f: y = 16'hfe00;
			16'ha280: y = 16'hfe00;
			16'ha281: y = 16'hfe00;
			16'ha282: y = 16'hfe00;
			16'ha283: y = 16'hfe00;
			16'ha284: y = 16'hfe00;
			16'ha285: y = 16'hfe00;
			16'ha286: y = 16'hfe00;
			16'ha287: y = 16'hfe00;
			16'ha288: y = 16'hfe00;
			16'ha289: y = 16'hfe00;
			16'ha28a: y = 16'hfe00;
			16'ha28b: y = 16'hfe00;
			16'ha28c: y = 16'hfe00;
			16'ha28d: y = 16'hfe00;
			16'ha28e: y = 16'hfe00;
			16'ha28f: y = 16'hfe00;
			16'ha290: y = 16'hfe00;
			16'ha291: y = 16'hfe00;
			16'ha292: y = 16'hfe00;
			16'ha293: y = 16'hfe00;
			16'ha294: y = 16'hfe00;
			16'ha295: y = 16'hfe00;
			16'ha296: y = 16'hfe00;
			16'ha297: y = 16'hfe00;
			16'ha298: y = 16'hfe00;
			16'ha299: y = 16'hfe00;
			16'ha29a: y = 16'hfe00;
			16'ha29b: y = 16'hfe00;
			16'ha29c: y = 16'hfe00;
			16'ha29d: y = 16'hfe00;
			16'ha29e: y = 16'hfe00;
			16'ha29f: y = 16'hfe00;
			16'ha2a0: y = 16'hfe00;
			16'ha2a1: y = 16'hfe00;
			16'ha2a2: y = 16'hfe00;
			16'ha2a3: y = 16'hfe00;
			16'ha2a4: y = 16'hfe00;
			16'ha2a5: y = 16'hfe00;
			16'ha2a6: y = 16'hfe00;
			16'ha2a7: y = 16'hfe00;
			16'ha2a8: y = 16'hfe00;
			16'ha2a9: y = 16'hfe00;
			16'ha2aa: y = 16'hfe00;
			16'ha2ab: y = 16'hfe00;
			16'ha2ac: y = 16'hfe00;
			16'ha2ad: y = 16'hfe00;
			16'ha2ae: y = 16'hfe00;
			16'ha2af: y = 16'hfe00;
			16'ha2b0: y = 16'hfe00;
			16'ha2b1: y = 16'hfe00;
			16'ha2b2: y = 16'hfe00;
			16'ha2b3: y = 16'hfe00;
			16'ha2b4: y = 16'hfe00;
			16'ha2b5: y = 16'hfe00;
			16'ha2b6: y = 16'hfe00;
			16'ha2b7: y = 16'hfe00;
			16'ha2b8: y = 16'hfe00;
			16'ha2b9: y = 16'hfe00;
			16'ha2ba: y = 16'hfe00;
			16'ha2bb: y = 16'hfe00;
			16'ha2bc: y = 16'hfe00;
			16'ha2bd: y = 16'hfe00;
			16'ha2be: y = 16'hfe00;
			16'ha2bf: y = 16'hfe00;
			16'ha2c0: y = 16'hfe00;
			16'ha2c1: y = 16'hfe00;
			16'ha2c2: y = 16'hfe00;
			16'ha2c3: y = 16'hfe00;
			16'ha2c4: y = 16'hfe00;
			16'ha2c5: y = 16'hfe00;
			16'ha2c6: y = 16'hfe00;
			16'ha2c7: y = 16'hfe00;
			16'ha2c8: y = 16'hfe00;
			16'ha2c9: y = 16'hfe00;
			16'ha2ca: y = 16'hfe00;
			16'ha2cb: y = 16'hfe00;
			16'ha2cc: y = 16'hfe00;
			16'ha2cd: y = 16'hfe00;
			16'ha2ce: y = 16'hfe00;
			16'ha2cf: y = 16'hfe00;
			16'ha2d0: y = 16'hfe00;
			16'ha2d1: y = 16'hfe00;
			16'ha2d2: y = 16'hfe00;
			16'ha2d3: y = 16'hfe00;
			16'ha2d4: y = 16'hfe00;
			16'ha2d5: y = 16'hfe00;
			16'ha2d6: y = 16'hfe00;
			16'ha2d7: y = 16'hfe00;
			16'ha2d8: y = 16'hfe00;
			16'ha2d9: y = 16'hfe00;
			16'ha2da: y = 16'hfe00;
			16'ha2db: y = 16'hfe00;
			16'ha2dc: y = 16'hfe00;
			16'ha2dd: y = 16'hfe00;
			16'ha2de: y = 16'hfe00;
			16'ha2df: y = 16'hfe00;
			16'ha2e0: y = 16'hfe00;
			16'ha2e1: y = 16'hfe00;
			16'ha2e2: y = 16'hfe00;
			16'ha2e3: y = 16'hfe00;
			16'ha2e4: y = 16'hfe00;
			16'ha2e5: y = 16'hfe00;
			16'ha2e6: y = 16'hfe00;
			16'ha2e7: y = 16'hfe00;
			16'ha2e8: y = 16'hfe00;
			16'ha2e9: y = 16'hfe00;
			16'ha2ea: y = 16'hfe00;
			16'ha2eb: y = 16'hfe00;
			16'ha2ec: y = 16'hfe00;
			16'ha2ed: y = 16'hfe00;
			16'ha2ee: y = 16'hfe00;
			16'ha2ef: y = 16'hfe00;
			16'ha2f0: y = 16'hfe00;
			16'ha2f1: y = 16'hfe00;
			16'ha2f2: y = 16'hfe00;
			16'ha2f3: y = 16'hfe00;
			16'ha2f4: y = 16'hfe00;
			16'ha2f5: y = 16'hfe00;
			16'ha2f6: y = 16'hfe00;
			16'ha2f7: y = 16'hfe00;
			16'ha2f8: y = 16'hfe00;
			16'ha2f9: y = 16'hfe00;
			16'ha2fa: y = 16'hfe00;
			16'ha2fb: y = 16'hfe00;
			16'ha2fc: y = 16'hfe00;
			16'ha2fd: y = 16'hfe00;
			16'ha2fe: y = 16'hfe00;
			16'ha2ff: y = 16'hfe00;
			16'ha300: y = 16'hfe00;
			16'ha301: y = 16'hfe00;
			16'ha302: y = 16'hfe00;
			16'ha303: y = 16'hfe00;
			16'ha304: y = 16'hfe00;
			16'ha305: y = 16'hfe00;
			16'ha306: y = 16'hfe00;
			16'ha307: y = 16'hfe00;
			16'ha308: y = 16'hfe00;
			16'ha309: y = 16'hfe00;
			16'ha30a: y = 16'hfe00;
			16'ha30b: y = 16'hfe00;
			16'ha30c: y = 16'hfe00;
			16'ha30d: y = 16'hfe00;
			16'ha30e: y = 16'hfe00;
			16'ha30f: y = 16'hfe00;
			16'ha310: y = 16'hfe00;
			16'ha311: y = 16'hfe00;
			16'ha312: y = 16'hfe00;
			16'ha313: y = 16'hfe00;
			16'ha314: y = 16'hfe00;
			16'ha315: y = 16'hfe00;
			16'ha316: y = 16'hfe00;
			16'ha317: y = 16'hfe00;
			16'ha318: y = 16'hfe00;
			16'ha319: y = 16'hfe00;
			16'ha31a: y = 16'hfe00;
			16'ha31b: y = 16'hfe00;
			16'ha31c: y = 16'hfe00;
			16'ha31d: y = 16'hfe00;
			16'ha31e: y = 16'hfe00;
			16'ha31f: y = 16'hfe00;
			16'ha320: y = 16'hfe00;
			16'ha321: y = 16'hfe00;
			16'ha322: y = 16'hfe00;
			16'ha323: y = 16'hfe00;
			16'ha324: y = 16'hfe00;
			16'ha325: y = 16'hfe00;
			16'ha326: y = 16'hfe00;
			16'ha327: y = 16'hfe00;
			16'ha328: y = 16'hfe00;
			16'ha329: y = 16'hfe00;
			16'ha32a: y = 16'hfe00;
			16'ha32b: y = 16'hfe00;
			16'ha32c: y = 16'hfe00;
			16'ha32d: y = 16'hfe00;
			16'ha32e: y = 16'hfe00;
			16'ha32f: y = 16'hfe00;
			16'ha330: y = 16'hfe00;
			16'ha331: y = 16'hfe00;
			16'ha332: y = 16'hfe00;
			16'ha333: y = 16'hfe00;
			16'ha334: y = 16'hfe00;
			16'ha335: y = 16'hfe00;
			16'ha336: y = 16'hfe00;
			16'ha337: y = 16'hfe00;
			16'ha338: y = 16'hfe00;
			16'ha339: y = 16'hfe00;
			16'ha33a: y = 16'hfe00;
			16'ha33b: y = 16'hfe00;
			16'ha33c: y = 16'hfe00;
			16'ha33d: y = 16'hfe00;
			16'ha33e: y = 16'hfe00;
			16'ha33f: y = 16'hfe00;
			16'ha340: y = 16'hfe00;
			16'ha341: y = 16'hfe00;
			16'ha342: y = 16'hfe00;
			16'ha343: y = 16'hfe00;
			16'ha344: y = 16'hfe00;
			16'ha345: y = 16'hfe00;
			16'ha346: y = 16'hfe00;
			16'ha347: y = 16'hfe00;
			16'ha348: y = 16'hfe00;
			16'ha349: y = 16'hfe00;
			16'ha34a: y = 16'hfe00;
			16'ha34b: y = 16'hfe00;
			16'ha34c: y = 16'hfe00;
			16'ha34d: y = 16'hfe00;
			16'ha34e: y = 16'hfe00;
			16'ha34f: y = 16'hfe00;
			16'ha350: y = 16'hfe00;
			16'ha351: y = 16'hfe00;
			16'ha352: y = 16'hfe00;
			16'ha353: y = 16'hfe00;
			16'ha354: y = 16'hfe00;
			16'ha355: y = 16'hfe00;
			16'ha356: y = 16'hfe00;
			16'ha357: y = 16'hfe00;
			16'ha358: y = 16'hfe00;
			16'ha359: y = 16'hfe00;
			16'ha35a: y = 16'hfe00;
			16'ha35b: y = 16'hfe00;
			16'ha35c: y = 16'hfe00;
			16'ha35d: y = 16'hfe00;
			16'ha35e: y = 16'hfe00;
			16'ha35f: y = 16'hfe00;
			16'ha360: y = 16'hfe00;
			16'ha361: y = 16'hfe00;
			16'ha362: y = 16'hfe00;
			16'ha363: y = 16'hfe00;
			16'ha364: y = 16'hfe00;
			16'ha365: y = 16'hfe00;
			16'ha366: y = 16'hfe00;
			16'ha367: y = 16'hfe00;
			16'ha368: y = 16'hfe00;
			16'ha369: y = 16'hfe00;
			16'ha36a: y = 16'hfe00;
			16'ha36b: y = 16'hfe00;
			16'ha36c: y = 16'hfe00;
			16'ha36d: y = 16'hfe00;
			16'ha36e: y = 16'hfe00;
			16'ha36f: y = 16'hfe00;
			16'ha370: y = 16'hfe00;
			16'ha371: y = 16'hfe00;
			16'ha372: y = 16'hfe00;
			16'ha373: y = 16'hfe00;
			16'ha374: y = 16'hfe00;
			16'ha375: y = 16'hfe00;
			16'ha376: y = 16'hfe00;
			16'ha377: y = 16'hfe00;
			16'ha378: y = 16'hfe00;
			16'ha379: y = 16'hfe00;
			16'ha37a: y = 16'hfe00;
			16'ha37b: y = 16'hfe00;
			16'ha37c: y = 16'hfe00;
			16'ha37d: y = 16'hfe00;
			16'ha37e: y = 16'hfe00;
			16'ha37f: y = 16'hfe00;
			16'ha380: y = 16'hfe00;
			16'ha381: y = 16'hfe00;
			16'ha382: y = 16'hfe00;
			16'ha383: y = 16'hfe00;
			16'ha384: y = 16'hfe00;
			16'ha385: y = 16'hfe00;
			16'ha386: y = 16'hfe00;
			16'ha387: y = 16'hfe00;
			16'ha388: y = 16'hfe00;
			16'ha389: y = 16'hfe00;
			16'ha38a: y = 16'hfe00;
			16'ha38b: y = 16'hfe00;
			16'ha38c: y = 16'hfe00;
			16'ha38d: y = 16'hfe00;
			16'ha38e: y = 16'hfe00;
			16'ha38f: y = 16'hfe00;
			16'ha390: y = 16'hfe00;
			16'ha391: y = 16'hfe00;
			16'ha392: y = 16'hfe00;
			16'ha393: y = 16'hfe00;
			16'ha394: y = 16'hfe00;
			16'ha395: y = 16'hfe00;
			16'ha396: y = 16'hfe00;
			16'ha397: y = 16'hfe00;
			16'ha398: y = 16'hfe00;
			16'ha399: y = 16'hfe00;
			16'ha39a: y = 16'hfe00;
			16'ha39b: y = 16'hfe00;
			16'ha39c: y = 16'hfe00;
			16'ha39d: y = 16'hfe00;
			16'ha39e: y = 16'hfe00;
			16'ha39f: y = 16'hfe00;
			16'ha3a0: y = 16'hfe00;
			16'ha3a1: y = 16'hfe00;
			16'ha3a2: y = 16'hfe00;
			16'ha3a3: y = 16'hfe00;
			16'ha3a4: y = 16'hfe00;
			16'ha3a5: y = 16'hfe00;
			16'ha3a6: y = 16'hfe00;
			16'ha3a7: y = 16'hfe00;
			16'ha3a8: y = 16'hfe00;
			16'ha3a9: y = 16'hfe00;
			16'ha3aa: y = 16'hfe00;
			16'ha3ab: y = 16'hfe00;
			16'ha3ac: y = 16'hfe00;
			16'ha3ad: y = 16'hfe00;
			16'ha3ae: y = 16'hfe00;
			16'ha3af: y = 16'hfe00;
			16'ha3b0: y = 16'hfe00;
			16'ha3b1: y = 16'hfe00;
			16'ha3b2: y = 16'hfe00;
			16'ha3b3: y = 16'hfe00;
			16'ha3b4: y = 16'hfe00;
			16'ha3b5: y = 16'hfe00;
			16'ha3b6: y = 16'hfe00;
			16'ha3b7: y = 16'hfe00;
			16'ha3b8: y = 16'hfe00;
			16'ha3b9: y = 16'hfe00;
			16'ha3ba: y = 16'hfe00;
			16'ha3bb: y = 16'hfe00;
			16'ha3bc: y = 16'hfe00;
			16'ha3bd: y = 16'hfe00;
			16'ha3be: y = 16'hfe00;
			16'ha3bf: y = 16'hfe00;
			16'ha3c0: y = 16'hfe00;
			16'ha3c1: y = 16'hfe00;
			16'ha3c2: y = 16'hfe00;
			16'ha3c3: y = 16'hfe00;
			16'ha3c4: y = 16'hfe00;
			16'ha3c5: y = 16'hfe00;
			16'ha3c6: y = 16'hfe00;
			16'ha3c7: y = 16'hfe00;
			16'ha3c8: y = 16'hfe00;
			16'ha3c9: y = 16'hfe00;
			16'ha3ca: y = 16'hfe00;
			16'ha3cb: y = 16'hfe00;
			16'ha3cc: y = 16'hfe00;
			16'ha3cd: y = 16'hfe00;
			16'ha3ce: y = 16'hfe00;
			16'ha3cf: y = 16'hfe00;
			16'ha3d0: y = 16'hfe00;
			16'ha3d1: y = 16'hfe00;
			16'ha3d2: y = 16'hfe00;
			16'ha3d3: y = 16'hfe00;
			16'ha3d4: y = 16'hfe00;
			16'ha3d5: y = 16'hfe00;
			16'ha3d6: y = 16'hfe00;
			16'ha3d7: y = 16'hfe00;
			16'ha3d8: y = 16'hfe00;
			16'ha3d9: y = 16'hfe00;
			16'ha3da: y = 16'hfe00;
			16'ha3db: y = 16'hfe00;
			16'ha3dc: y = 16'hfe00;
			16'ha3dd: y = 16'hfe00;
			16'ha3de: y = 16'hfe00;
			16'ha3df: y = 16'hfe00;
			16'ha3e0: y = 16'hfe00;
			16'ha3e1: y = 16'hfe00;
			16'ha3e2: y = 16'hfe00;
			16'ha3e3: y = 16'hfe00;
			16'ha3e4: y = 16'hfe00;
			16'ha3e5: y = 16'hfe00;
			16'ha3e6: y = 16'hfe00;
			16'ha3e7: y = 16'hfe00;
			16'ha3e8: y = 16'hfe00;
			16'ha3e9: y = 16'hfe00;
			16'ha3ea: y = 16'hfe00;
			16'ha3eb: y = 16'hfe00;
			16'ha3ec: y = 16'hfe00;
			16'ha3ed: y = 16'hfe00;
			16'ha3ee: y = 16'hfe00;
			16'ha3ef: y = 16'hfe00;
			16'ha3f0: y = 16'hfe00;
			16'ha3f1: y = 16'hfe00;
			16'ha3f2: y = 16'hfe00;
			16'ha3f3: y = 16'hfe00;
			16'ha3f4: y = 16'hfe00;
			16'ha3f5: y = 16'hfe00;
			16'ha3f6: y = 16'hfe00;
			16'ha3f7: y = 16'hfe00;
			16'ha3f8: y = 16'hfe00;
			16'ha3f9: y = 16'hfe00;
			16'ha3fa: y = 16'hfe00;
			16'ha3fb: y = 16'hfe00;
			16'ha3fc: y = 16'hfe00;
			16'ha3fd: y = 16'hfe00;
			16'ha3fe: y = 16'hfe00;
			16'ha3ff: y = 16'hfe00;
			16'ha400: y = 16'hfe00;
			16'ha401: y = 16'hfe00;
			16'ha402: y = 16'hfe00;
			16'ha403: y = 16'hfe00;
			16'ha404: y = 16'hfe00;
			16'ha405: y = 16'hfe00;
			16'ha406: y = 16'hfe00;
			16'ha407: y = 16'hfe00;
			16'ha408: y = 16'hfe00;
			16'ha409: y = 16'hfe00;
			16'ha40a: y = 16'hfe00;
			16'ha40b: y = 16'hfe00;
			16'ha40c: y = 16'hfe00;
			16'ha40d: y = 16'hfe00;
			16'ha40e: y = 16'hfe00;
			16'ha40f: y = 16'hfe00;
			16'ha410: y = 16'hfe00;
			16'ha411: y = 16'hfe00;
			16'ha412: y = 16'hfe00;
			16'ha413: y = 16'hfe00;
			16'ha414: y = 16'hfe00;
			16'ha415: y = 16'hfe00;
			16'ha416: y = 16'hfe00;
			16'ha417: y = 16'hfe00;
			16'ha418: y = 16'hfe00;
			16'ha419: y = 16'hfe00;
			16'ha41a: y = 16'hfe00;
			16'ha41b: y = 16'hfe00;
			16'ha41c: y = 16'hfe00;
			16'ha41d: y = 16'hfe00;
			16'ha41e: y = 16'hfe00;
			16'ha41f: y = 16'hfe00;
			16'ha420: y = 16'hfe00;
			16'ha421: y = 16'hfe00;
			16'ha422: y = 16'hfe00;
			16'ha423: y = 16'hfe00;
			16'ha424: y = 16'hfe00;
			16'ha425: y = 16'hfe00;
			16'ha426: y = 16'hfe00;
			16'ha427: y = 16'hfe00;
			16'ha428: y = 16'hfe00;
			16'ha429: y = 16'hfe00;
			16'ha42a: y = 16'hfe00;
			16'ha42b: y = 16'hfe00;
			16'ha42c: y = 16'hfe00;
			16'ha42d: y = 16'hfe00;
			16'ha42e: y = 16'hfe00;
			16'ha42f: y = 16'hfe00;
			16'ha430: y = 16'hfe00;
			16'ha431: y = 16'hfe00;
			16'ha432: y = 16'hfe00;
			16'ha433: y = 16'hfe00;
			16'ha434: y = 16'hfe00;
			16'ha435: y = 16'hfe00;
			16'ha436: y = 16'hfe00;
			16'ha437: y = 16'hfe00;
			16'ha438: y = 16'hfe00;
			16'ha439: y = 16'hfe00;
			16'ha43a: y = 16'hfe00;
			16'ha43b: y = 16'hfe00;
			16'ha43c: y = 16'hfe00;
			16'ha43d: y = 16'hfe00;
			16'ha43e: y = 16'hfe00;
			16'ha43f: y = 16'hfe00;
			16'ha440: y = 16'hfe00;
			16'ha441: y = 16'hfe00;
			16'ha442: y = 16'hfe00;
			16'ha443: y = 16'hfe00;
			16'ha444: y = 16'hfe00;
			16'ha445: y = 16'hfe00;
			16'ha446: y = 16'hfe00;
			16'ha447: y = 16'hfe00;
			16'ha448: y = 16'hfe00;
			16'ha449: y = 16'hfe00;
			16'ha44a: y = 16'hfe00;
			16'ha44b: y = 16'hfe00;
			16'ha44c: y = 16'hfe00;
			16'ha44d: y = 16'hfe00;
			16'ha44e: y = 16'hfe00;
			16'ha44f: y = 16'hfe00;
			16'ha450: y = 16'hfe00;
			16'ha451: y = 16'hfe00;
			16'ha452: y = 16'hfe00;
			16'ha453: y = 16'hfe00;
			16'ha454: y = 16'hfe00;
			16'ha455: y = 16'hfe00;
			16'ha456: y = 16'hfe00;
			16'ha457: y = 16'hfe00;
			16'ha458: y = 16'hfe00;
			16'ha459: y = 16'hfe00;
			16'ha45a: y = 16'hfe00;
			16'ha45b: y = 16'hfe00;
			16'ha45c: y = 16'hfe00;
			16'ha45d: y = 16'hfe00;
			16'ha45e: y = 16'hfe00;
			16'ha45f: y = 16'hfe00;
			16'ha460: y = 16'hfe00;
			16'ha461: y = 16'hfe00;
			16'ha462: y = 16'hfe00;
			16'ha463: y = 16'hfe00;
			16'ha464: y = 16'hfe00;
			16'ha465: y = 16'hfe00;
			16'ha466: y = 16'hfe00;
			16'ha467: y = 16'hfe00;
			16'ha468: y = 16'hfe00;
			16'ha469: y = 16'hfe00;
			16'ha46a: y = 16'hfe00;
			16'ha46b: y = 16'hfe00;
			16'ha46c: y = 16'hfe00;
			16'ha46d: y = 16'hfe00;
			16'ha46e: y = 16'hfe00;
			16'ha46f: y = 16'hfe00;
			16'ha470: y = 16'hfe00;
			16'ha471: y = 16'hfe00;
			16'ha472: y = 16'hfe00;
			16'ha473: y = 16'hfe00;
			16'ha474: y = 16'hfe00;
			16'ha475: y = 16'hfe00;
			16'ha476: y = 16'hfe00;
			16'ha477: y = 16'hfe00;
			16'ha478: y = 16'hfe00;
			16'ha479: y = 16'hfe00;
			16'ha47a: y = 16'hfe00;
			16'ha47b: y = 16'hfe00;
			16'ha47c: y = 16'hfe00;
			16'ha47d: y = 16'hfe00;
			16'ha47e: y = 16'hfe00;
			16'ha47f: y = 16'hfe00;
			16'ha480: y = 16'hfe00;
			16'ha481: y = 16'hfe00;
			16'ha482: y = 16'hfe00;
			16'ha483: y = 16'hfe00;
			16'ha484: y = 16'hfe00;
			16'ha485: y = 16'hfe00;
			16'ha486: y = 16'hfe00;
			16'ha487: y = 16'hfe00;
			16'ha488: y = 16'hfe00;
			16'ha489: y = 16'hfe00;
			16'ha48a: y = 16'hfe00;
			16'ha48b: y = 16'hfe00;
			16'ha48c: y = 16'hfe00;
			16'ha48d: y = 16'hfe00;
			16'ha48e: y = 16'hfe00;
			16'ha48f: y = 16'hfe00;
			16'ha490: y = 16'hfe00;
			16'ha491: y = 16'hfe00;
			16'ha492: y = 16'hfe00;
			16'ha493: y = 16'hfe00;
			16'ha494: y = 16'hfe00;
			16'ha495: y = 16'hfe00;
			16'ha496: y = 16'hfe00;
			16'ha497: y = 16'hfe00;
			16'ha498: y = 16'hfe00;
			16'ha499: y = 16'hfe00;
			16'ha49a: y = 16'hfe00;
			16'ha49b: y = 16'hfe00;
			16'ha49c: y = 16'hfe00;
			16'ha49d: y = 16'hfe00;
			16'ha49e: y = 16'hfe00;
			16'ha49f: y = 16'hfe00;
			16'ha4a0: y = 16'hfe00;
			16'ha4a1: y = 16'hfe00;
			16'ha4a2: y = 16'hfe00;
			16'ha4a3: y = 16'hfe00;
			16'ha4a4: y = 16'hfe00;
			16'ha4a5: y = 16'hfe00;
			16'ha4a6: y = 16'hfe00;
			16'ha4a7: y = 16'hfe00;
			16'ha4a8: y = 16'hfe00;
			16'ha4a9: y = 16'hfe00;
			16'ha4aa: y = 16'hfe00;
			16'ha4ab: y = 16'hfe00;
			16'ha4ac: y = 16'hfe00;
			16'ha4ad: y = 16'hfe00;
			16'ha4ae: y = 16'hfe00;
			16'ha4af: y = 16'hfe00;
			16'ha4b0: y = 16'hfe00;
			16'ha4b1: y = 16'hfe00;
			16'ha4b2: y = 16'hfe00;
			16'ha4b3: y = 16'hfe00;
			16'ha4b4: y = 16'hfe00;
			16'ha4b5: y = 16'hfe00;
			16'ha4b6: y = 16'hfe00;
			16'ha4b7: y = 16'hfe00;
			16'ha4b8: y = 16'hfe00;
			16'ha4b9: y = 16'hfe00;
			16'ha4ba: y = 16'hfe00;
			16'ha4bb: y = 16'hfe00;
			16'ha4bc: y = 16'hfe00;
			16'ha4bd: y = 16'hfe00;
			16'ha4be: y = 16'hfe00;
			16'ha4bf: y = 16'hfe00;
			16'ha4c0: y = 16'hfe00;
			16'ha4c1: y = 16'hfe00;
			16'ha4c2: y = 16'hfe00;
			16'ha4c3: y = 16'hfe00;
			16'ha4c4: y = 16'hfe00;
			16'ha4c5: y = 16'hfe00;
			16'ha4c6: y = 16'hfe00;
			16'ha4c7: y = 16'hfe00;
			16'ha4c8: y = 16'hfe00;
			16'ha4c9: y = 16'hfe00;
			16'ha4ca: y = 16'hfe00;
			16'ha4cb: y = 16'hfe00;
			16'ha4cc: y = 16'hfe00;
			16'ha4cd: y = 16'hfe00;
			16'ha4ce: y = 16'hfe00;
			16'ha4cf: y = 16'hfe00;
			16'ha4d0: y = 16'hfe00;
			16'ha4d1: y = 16'hfe00;
			16'ha4d2: y = 16'hfe00;
			16'ha4d3: y = 16'hfe00;
			16'ha4d4: y = 16'hfe00;
			16'ha4d5: y = 16'hfe00;
			16'ha4d6: y = 16'hfe00;
			16'ha4d7: y = 16'hfe00;
			16'ha4d8: y = 16'hfe00;
			16'ha4d9: y = 16'hfe00;
			16'ha4da: y = 16'hfe00;
			16'ha4db: y = 16'hfe00;
			16'ha4dc: y = 16'hfe00;
			16'ha4dd: y = 16'hfe00;
			16'ha4de: y = 16'hfe00;
			16'ha4df: y = 16'hfe00;
			16'ha4e0: y = 16'hfe00;
			16'ha4e1: y = 16'hfe00;
			16'ha4e2: y = 16'hfe00;
			16'ha4e3: y = 16'hfe00;
			16'ha4e4: y = 16'hfe00;
			16'ha4e5: y = 16'hfe00;
			16'ha4e6: y = 16'hfe00;
			16'ha4e7: y = 16'hfe00;
			16'ha4e8: y = 16'hfe00;
			16'ha4e9: y = 16'hfe00;
			16'ha4ea: y = 16'hfe00;
			16'ha4eb: y = 16'hfe00;
			16'ha4ec: y = 16'hfe00;
			16'ha4ed: y = 16'hfe00;
			16'ha4ee: y = 16'hfe00;
			16'ha4ef: y = 16'hfe00;
			16'ha4f0: y = 16'hfe00;
			16'ha4f1: y = 16'hfe00;
			16'ha4f2: y = 16'hfe00;
			16'ha4f3: y = 16'hfe00;
			16'ha4f4: y = 16'hfe00;
			16'ha4f5: y = 16'hfe00;
			16'ha4f6: y = 16'hfe00;
			16'ha4f7: y = 16'hfe00;
			16'ha4f8: y = 16'hfe00;
			16'ha4f9: y = 16'hfe00;
			16'ha4fa: y = 16'hfe00;
			16'ha4fb: y = 16'hfe00;
			16'ha4fc: y = 16'hfe00;
			16'ha4fd: y = 16'hfe00;
			16'ha4fe: y = 16'hfe00;
			16'ha4ff: y = 16'hfe00;
			16'ha500: y = 16'hfe00;
			16'ha501: y = 16'hfe00;
			16'ha502: y = 16'hfe00;
			16'ha503: y = 16'hfe00;
			16'ha504: y = 16'hfe00;
			16'ha505: y = 16'hfe00;
			16'ha506: y = 16'hfe00;
			16'ha507: y = 16'hfe00;
			16'ha508: y = 16'hfe00;
			16'ha509: y = 16'hfe00;
			16'ha50a: y = 16'hfe00;
			16'ha50b: y = 16'hfe00;
			16'ha50c: y = 16'hfe00;
			16'ha50d: y = 16'hfe00;
			16'ha50e: y = 16'hfe00;
			16'ha50f: y = 16'hfe00;
			16'ha510: y = 16'hfe00;
			16'ha511: y = 16'hfe00;
			16'ha512: y = 16'hfe00;
			16'ha513: y = 16'hfe00;
			16'ha514: y = 16'hfe00;
			16'ha515: y = 16'hfe00;
			16'ha516: y = 16'hfe00;
			16'ha517: y = 16'hfe00;
			16'ha518: y = 16'hfe00;
			16'ha519: y = 16'hfe00;
			16'ha51a: y = 16'hfe00;
			16'ha51b: y = 16'hfe00;
			16'ha51c: y = 16'hfe00;
			16'ha51d: y = 16'hfe00;
			16'ha51e: y = 16'hfe00;
			16'ha51f: y = 16'hfe00;
			16'ha520: y = 16'hfe00;
			16'ha521: y = 16'hfe00;
			16'ha522: y = 16'hfe00;
			16'ha523: y = 16'hfe00;
			16'ha524: y = 16'hfe00;
			16'ha525: y = 16'hfe00;
			16'ha526: y = 16'hfe00;
			16'ha527: y = 16'hfe00;
			16'ha528: y = 16'hfe00;
			16'ha529: y = 16'hfe00;
			16'ha52a: y = 16'hfe00;
			16'ha52b: y = 16'hfe00;
			16'ha52c: y = 16'hfe00;
			16'ha52d: y = 16'hfe00;
			16'ha52e: y = 16'hfe00;
			16'ha52f: y = 16'hfe00;
			16'ha530: y = 16'hfe00;
			16'ha531: y = 16'hfe00;
			16'ha532: y = 16'hfe00;
			16'ha533: y = 16'hfe00;
			16'ha534: y = 16'hfe00;
			16'ha535: y = 16'hfe00;
			16'ha536: y = 16'hfe00;
			16'ha537: y = 16'hfe00;
			16'ha538: y = 16'hfe00;
			16'ha539: y = 16'hfe00;
			16'ha53a: y = 16'hfe00;
			16'ha53b: y = 16'hfe00;
			16'ha53c: y = 16'hfe00;
			16'ha53d: y = 16'hfe00;
			16'ha53e: y = 16'hfe00;
			16'ha53f: y = 16'hfe00;
			16'ha540: y = 16'hfe00;
			16'ha541: y = 16'hfe00;
			16'ha542: y = 16'hfe00;
			16'ha543: y = 16'hfe00;
			16'ha544: y = 16'hfe00;
			16'ha545: y = 16'hfe00;
			16'ha546: y = 16'hfe00;
			16'ha547: y = 16'hfe00;
			16'ha548: y = 16'hfe00;
			16'ha549: y = 16'hfe00;
			16'ha54a: y = 16'hfe00;
			16'ha54b: y = 16'hfe00;
			16'ha54c: y = 16'hfe00;
			16'ha54d: y = 16'hfe00;
			16'ha54e: y = 16'hfe00;
			16'ha54f: y = 16'hfe00;
			16'ha550: y = 16'hfe00;
			16'ha551: y = 16'hfe00;
			16'ha552: y = 16'hfe00;
			16'ha553: y = 16'hfe00;
			16'ha554: y = 16'hfe00;
			16'ha555: y = 16'hfe00;
			16'ha556: y = 16'hfe00;
			16'ha557: y = 16'hfe00;
			16'ha558: y = 16'hfe00;
			16'ha559: y = 16'hfe00;
			16'ha55a: y = 16'hfe00;
			16'ha55b: y = 16'hfe00;
			16'ha55c: y = 16'hfe00;
			16'ha55d: y = 16'hfe00;
			16'ha55e: y = 16'hfe00;
			16'ha55f: y = 16'hfe00;
			16'ha560: y = 16'hfe00;
			16'ha561: y = 16'hfe00;
			16'ha562: y = 16'hfe00;
			16'ha563: y = 16'hfe00;
			16'ha564: y = 16'hfe00;
			16'ha565: y = 16'hfe00;
			16'ha566: y = 16'hfe00;
			16'ha567: y = 16'hfe00;
			16'ha568: y = 16'hfe00;
			16'ha569: y = 16'hfe00;
			16'ha56a: y = 16'hfe00;
			16'ha56b: y = 16'hfe00;
			16'ha56c: y = 16'hfe00;
			16'ha56d: y = 16'hfe00;
			16'ha56e: y = 16'hfe00;
			16'ha56f: y = 16'hfe00;
			16'ha570: y = 16'hfe00;
			16'ha571: y = 16'hfe00;
			16'ha572: y = 16'hfe00;
			16'ha573: y = 16'hfe00;
			16'ha574: y = 16'hfe00;
			16'ha575: y = 16'hfe00;
			16'ha576: y = 16'hfe00;
			16'ha577: y = 16'hfe00;
			16'ha578: y = 16'hfe00;
			16'ha579: y = 16'hfe00;
			16'ha57a: y = 16'hfe00;
			16'ha57b: y = 16'hfe00;
			16'ha57c: y = 16'hfe00;
			16'ha57d: y = 16'hfe00;
			16'ha57e: y = 16'hfe00;
			16'ha57f: y = 16'hfe00;
			16'ha580: y = 16'hfe00;
			16'ha581: y = 16'hfe00;
			16'ha582: y = 16'hfe00;
			16'ha583: y = 16'hfe00;
			16'ha584: y = 16'hfe00;
			16'ha585: y = 16'hfe00;
			16'ha586: y = 16'hfe00;
			16'ha587: y = 16'hfe00;
			16'ha588: y = 16'hfe00;
			16'ha589: y = 16'hfe00;
			16'ha58a: y = 16'hfe00;
			16'ha58b: y = 16'hfe00;
			16'ha58c: y = 16'hfe00;
			16'ha58d: y = 16'hfe00;
			16'ha58e: y = 16'hfe00;
			16'ha58f: y = 16'hfe00;
			16'ha590: y = 16'hfe00;
			16'ha591: y = 16'hfe00;
			16'ha592: y = 16'hfe00;
			16'ha593: y = 16'hfe00;
			16'ha594: y = 16'hfe00;
			16'ha595: y = 16'hfe00;
			16'ha596: y = 16'hfe00;
			16'ha597: y = 16'hfe00;
			16'ha598: y = 16'hfe00;
			16'ha599: y = 16'hfe00;
			16'ha59a: y = 16'hfe00;
			16'ha59b: y = 16'hfe00;
			16'ha59c: y = 16'hfe00;
			16'ha59d: y = 16'hfe00;
			16'ha59e: y = 16'hfe00;
			16'ha59f: y = 16'hfe00;
			16'ha5a0: y = 16'hfe00;
			16'ha5a1: y = 16'hfe00;
			16'ha5a2: y = 16'hfe00;
			16'ha5a3: y = 16'hfe00;
			16'ha5a4: y = 16'hfe00;
			16'ha5a5: y = 16'hfe00;
			16'ha5a6: y = 16'hfe00;
			16'ha5a7: y = 16'hfe00;
			16'ha5a8: y = 16'hfe00;
			16'ha5a9: y = 16'hfe00;
			16'ha5aa: y = 16'hfe00;
			16'ha5ab: y = 16'hfe00;
			16'ha5ac: y = 16'hfe00;
			16'ha5ad: y = 16'hfe00;
			16'ha5ae: y = 16'hfe00;
			16'ha5af: y = 16'hfe00;
			16'ha5b0: y = 16'hfe00;
			16'ha5b1: y = 16'hfe00;
			16'ha5b2: y = 16'hfe00;
			16'ha5b3: y = 16'hfe00;
			16'ha5b4: y = 16'hfe00;
			16'ha5b5: y = 16'hfe00;
			16'ha5b6: y = 16'hfe00;
			16'ha5b7: y = 16'hfe00;
			16'ha5b8: y = 16'hfe00;
			16'ha5b9: y = 16'hfe00;
			16'ha5ba: y = 16'hfe00;
			16'ha5bb: y = 16'hfe00;
			16'ha5bc: y = 16'hfe00;
			16'ha5bd: y = 16'hfe00;
			16'ha5be: y = 16'hfe00;
			16'ha5bf: y = 16'hfe00;
			16'ha5c0: y = 16'hfe00;
			16'ha5c1: y = 16'hfe00;
			16'ha5c2: y = 16'hfe00;
			16'ha5c3: y = 16'hfe00;
			16'ha5c4: y = 16'hfe00;
			16'ha5c5: y = 16'hfe00;
			16'ha5c6: y = 16'hfe00;
			16'ha5c7: y = 16'hfe00;
			16'ha5c8: y = 16'hfe00;
			16'ha5c9: y = 16'hfe00;
			16'ha5ca: y = 16'hfe00;
			16'ha5cb: y = 16'hfe00;
			16'ha5cc: y = 16'hfe00;
			16'ha5cd: y = 16'hfe00;
			16'ha5ce: y = 16'hfe00;
			16'ha5cf: y = 16'hfe00;
			16'ha5d0: y = 16'hfe00;
			16'ha5d1: y = 16'hfe00;
			16'ha5d2: y = 16'hfe00;
			16'ha5d3: y = 16'hfe00;
			16'ha5d4: y = 16'hfe00;
			16'ha5d5: y = 16'hfe00;
			16'ha5d6: y = 16'hfe00;
			16'ha5d7: y = 16'hfe00;
			16'ha5d8: y = 16'hfe00;
			16'ha5d9: y = 16'hfe00;
			16'ha5da: y = 16'hfe00;
			16'ha5db: y = 16'hfe00;
			16'ha5dc: y = 16'hfe00;
			16'ha5dd: y = 16'hfe00;
			16'ha5de: y = 16'hfe00;
			16'ha5df: y = 16'hfe00;
			16'ha5e0: y = 16'hfe00;
			16'ha5e1: y = 16'hfe00;
			16'ha5e2: y = 16'hfe00;
			16'ha5e3: y = 16'hfe00;
			16'ha5e4: y = 16'hfe00;
			16'ha5e5: y = 16'hfe00;
			16'ha5e6: y = 16'hfe00;
			16'ha5e7: y = 16'hfe00;
			16'ha5e8: y = 16'hfe00;
			16'ha5e9: y = 16'hfe00;
			16'ha5ea: y = 16'hfe00;
			16'ha5eb: y = 16'hfe00;
			16'ha5ec: y = 16'hfe00;
			16'ha5ed: y = 16'hfe00;
			16'ha5ee: y = 16'hfe00;
			16'ha5ef: y = 16'hfe00;
			16'ha5f0: y = 16'hfe00;
			16'ha5f1: y = 16'hfe00;
			16'ha5f2: y = 16'hfe00;
			16'ha5f3: y = 16'hfe00;
			16'ha5f4: y = 16'hfe00;
			16'ha5f5: y = 16'hfe00;
			16'ha5f6: y = 16'hfe00;
			16'ha5f7: y = 16'hfe00;
			16'ha5f8: y = 16'hfe00;
			16'ha5f9: y = 16'hfe00;
			16'ha5fa: y = 16'hfe00;
			16'ha5fb: y = 16'hfe00;
			16'ha5fc: y = 16'hfe00;
			16'ha5fd: y = 16'hfe00;
			16'ha5fe: y = 16'hfe00;
			16'ha5ff: y = 16'hfe00;
			16'ha600: y = 16'hfe00;
			16'ha601: y = 16'hfe00;
			16'ha602: y = 16'hfe00;
			16'ha603: y = 16'hfe00;
			16'ha604: y = 16'hfe00;
			16'ha605: y = 16'hfe00;
			16'ha606: y = 16'hfe00;
			16'ha607: y = 16'hfe00;
			16'ha608: y = 16'hfe00;
			16'ha609: y = 16'hfe00;
			16'ha60a: y = 16'hfe00;
			16'ha60b: y = 16'hfe00;
			16'ha60c: y = 16'hfe00;
			16'ha60d: y = 16'hfe00;
			16'ha60e: y = 16'hfe00;
			16'ha60f: y = 16'hfe00;
			16'ha610: y = 16'hfe00;
			16'ha611: y = 16'hfe00;
			16'ha612: y = 16'hfe00;
			16'ha613: y = 16'hfe00;
			16'ha614: y = 16'hfe00;
			16'ha615: y = 16'hfe00;
			16'ha616: y = 16'hfe00;
			16'ha617: y = 16'hfe00;
			16'ha618: y = 16'hfe00;
			16'ha619: y = 16'hfe00;
			16'ha61a: y = 16'hfe00;
			16'ha61b: y = 16'hfe00;
			16'ha61c: y = 16'hfe00;
			16'ha61d: y = 16'hfe00;
			16'ha61e: y = 16'hfe00;
			16'ha61f: y = 16'hfe00;
			16'ha620: y = 16'hfe00;
			16'ha621: y = 16'hfe00;
			16'ha622: y = 16'hfe00;
			16'ha623: y = 16'hfe00;
			16'ha624: y = 16'hfe00;
			16'ha625: y = 16'hfe00;
			16'ha626: y = 16'hfe00;
			16'ha627: y = 16'hfe00;
			16'ha628: y = 16'hfe00;
			16'ha629: y = 16'hfe00;
			16'ha62a: y = 16'hfe00;
			16'ha62b: y = 16'hfe00;
			16'ha62c: y = 16'hfe00;
			16'ha62d: y = 16'hfe00;
			16'ha62e: y = 16'hfe00;
			16'ha62f: y = 16'hfe00;
			16'ha630: y = 16'hfe00;
			16'ha631: y = 16'hfe00;
			16'ha632: y = 16'hfe00;
			16'ha633: y = 16'hfe00;
			16'ha634: y = 16'hfe00;
			16'ha635: y = 16'hfe00;
			16'ha636: y = 16'hfe00;
			16'ha637: y = 16'hfe00;
			16'ha638: y = 16'hfe00;
			16'ha639: y = 16'hfe00;
			16'ha63a: y = 16'hfe00;
			16'ha63b: y = 16'hfe00;
			16'ha63c: y = 16'hfe00;
			16'ha63d: y = 16'hfe00;
			16'ha63e: y = 16'hfe00;
			16'ha63f: y = 16'hfe00;
			16'ha640: y = 16'hfe00;
			16'ha641: y = 16'hfe00;
			16'ha642: y = 16'hfe00;
			16'ha643: y = 16'hfe00;
			16'ha644: y = 16'hfe00;
			16'ha645: y = 16'hfe00;
			16'ha646: y = 16'hfe00;
			16'ha647: y = 16'hfe00;
			16'ha648: y = 16'hfe00;
			16'ha649: y = 16'hfe00;
			16'ha64a: y = 16'hfe00;
			16'ha64b: y = 16'hfe00;
			16'ha64c: y = 16'hfe00;
			16'ha64d: y = 16'hfe00;
			16'ha64e: y = 16'hfe00;
			16'ha64f: y = 16'hfe00;
			16'ha650: y = 16'hfe00;
			16'ha651: y = 16'hfe00;
			16'ha652: y = 16'hfe00;
			16'ha653: y = 16'hfe00;
			16'ha654: y = 16'hfe00;
			16'ha655: y = 16'hfe00;
			16'ha656: y = 16'hfe00;
			16'ha657: y = 16'hfe00;
			16'ha658: y = 16'hfe00;
			16'ha659: y = 16'hfe00;
			16'ha65a: y = 16'hfe00;
			16'ha65b: y = 16'hfe00;
			16'ha65c: y = 16'hfe00;
			16'ha65d: y = 16'hfe00;
			16'ha65e: y = 16'hfe00;
			16'ha65f: y = 16'hfe00;
			16'ha660: y = 16'hfe00;
			16'ha661: y = 16'hfe00;
			16'ha662: y = 16'hfe00;
			16'ha663: y = 16'hfe00;
			16'ha664: y = 16'hfe00;
			16'ha665: y = 16'hfe00;
			16'ha666: y = 16'hfe00;
			16'ha667: y = 16'hfe00;
			16'ha668: y = 16'hfe00;
			16'ha669: y = 16'hfe00;
			16'ha66a: y = 16'hfe00;
			16'ha66b: y = 16'hfe00;
			16'ha66c: y = 16'hfe00;
			16'ha66d: y = 16'hfe00;
			16'ha66e: y = 16'hfe00;
			16'ha66f: y = 16'hfe00;
			16'ha670: y = 16'hfe00;
			16'ha671: y = 16'hfe00;
			16'ha672: y = 16'hfe00;
			16'ha673: y = 16'hfe00;
			16'ha674: y = 16'hfe00;
			16'ha675: y = 16'hfe00;
			16'ha676: y = 16'hfe00;
			16'ha677: y = 16'hfe00;
			16'ha678: y = 16'hfe00;
			16'ha679: y = 16'hfe00;
			16'ha67a: y = 16'hfe00;
			16'ha67b: y = 16'hfe00;
			16'ha67c: y = 16'hfe00;
			16'ha67d: y = 16'hfe00;
			16'ha67e: y = 16'hfe00;
			16'ha67f: y = 16'hfe00;
			16'ha680: y = 16'hfe00;
			16'ha681: y = 16'hfe00;
			16'ha682: y = 16'hfe00;
			16'ha683: y = 16'hfe00;
			16'ha684: y = 16'hfe00;
			16'ha685: y = 16'hfe00;
			16'ha686: y = 16'hfe00;
			16'ha687: y = 16'hfe00;
			16'ha688: y = 16'hfe00;
			16'ha689: y = 16'hfe00;
			16'ha68a: y = 16'hfe00;
			16'ha68b: y = 16'hfe00;
			16'ha68c: y = 16'hfe00;
			16'ha68d: y = 16'hfe00;
			16'ha68e: y = 16'hfe00;
			16'ha68f: y = 16'hfe00;
			16'ha690: y = 16'hfe00;
			16'ha691: y = 16'hfe00;
			16'ha692: y = 16'hfe00;
			16'ha693: y = 16'hfe00;
			16'ha694: y = 16'hfe00;
			16'ha695: y = 16'hfe00;
			16'ha696: y = 16'hfe00;
			16'ha697: y = 16'hfe00;
			16'ha698: y = 16'hfe00;
			16'ha699: y = 16'hfe00;
			16'ha69a: y = 16'hfe00;
			16'ha69b: y = 16'hfe00;
			16'ha69c: y = 16'hfe00;
			16'ha69d: y = 16'hfe00;
			16'ha69e: y = 16'hfe00;
			16'ha69f: y = 16'hfe00;
			16'ha6a0: y = 16'hfe00;
			16'ha6a1: y = 16'hfe00;
			16'ha6a2: y = 16'hfe00;
			16'ha6a3: y = 16'hfe00;
			16'ha6a4: y = 16'hfe00;
			16'ha6a5: y = 16'hfe00;
			16'ha6a6: y = 16'hfe00;
			16'ha6a7: y = 16'hfe00;
			16'ha6a8: y = 16'hfe00;
			16'ha6a9: y = 16'hfe00;
			16'ha6aa: y = 16'hfe00;
			16'ha6ab: y = 16'hfe00;
			16'ha6ac: y = 16'hfe00;
			16'ha6ad: y = 16'hfe00;
			16'ha6ae: y = 16'hfe00;
			16'ha6af: y = 16'hfe00;
			16'ha6b0: y = 16'hfe00;
			16'ha6b1: y = 16'hfe00;
			16'ha6b2: y = 16'hfe00;
			16'ha6b3: y = 16'hfe00;
			16'ha6b4: y = 16'hfe00;
			16'ha6b5: y = 16'hfe00;
			16'ha6b6: y = 16'hfe00;
			16'ha6b7: y = 16'hfe00;
			16'ha6b8: y = 16'hfe00;
			16'ha6b9: y = 16'hfe00;
			16'ha6ba: y = 16'hfe00;
			16'ha6bb: y = 16'hfe00;
			16'ha6bc: y = 16'hfe00;
			16'ha6bd: y = 16'hfe00;
			16'ha6be: y = 16'hfe00;
			16'ha6bf: y = 16'hfe00;
			16'ha6c0: y = 16'hfe00;
			16'ha6c1: y = 16'hfe00;
			16'ha6c2: y = 16'hfe00;
			16'ha6c3: y = 16'hfe00;
			16'ha6c4: y = 16'hfe00;
			16'ha6c5: y = 16'hfe00;
			16'ha6c6: y = 16'hfe00;
			16'ha6c7: y = 16'hfe00;
			16'ha6c8: y = 16'hfe00;
			16'ha6c9: y = 16'hfe00;
			16'ha6ca: y = 16'hfe00;
			16'ha6cb: y = 16'hfe00;
			16'ha6cc: y = 16'hfe00;
			16'ha6cd: y = 16'hfe00;
			16'ha6ce: y = 16'hfe00;
			16'ha6cf: y = 16'hfe00;
			16'ha6d0: y = 16'hfe00;
			16'ha6d1: y = 16'hfe00;
			16'ha6d2: y = 16'hfe00;
			16'ha6d3: y = 16'hfe00;
			16'ha6d4: y = 16'hfe00;
			16'ha6d5: y = 16'hfe00;
			16'ha6d6: y = 16'hfe00;
			16'ha6d7: y = 16'hfe00;
			16'ha6d8: y = 16'hfe00;
			16'ha6d9: y = 16'hfe00;
			16'ha6da: y = 16'hfe00;
			16'ha6db: y = 16'hfe00;
			16'ha6dc: y = 16'hfe00;
			16'ha6dd: y = 16'hfe00;
			16'ha6de: y = 16'hfe00;
			16'ha6df: y = 16'hfe00;
			16'ha6e0: y = 16'hfe00;
			16'ha6e1: y = 16'hfe00;
			16'ha6e2: y = 16'hfe00;
			16'ha6e3: y = 16'hfe00;
			16'ha6e4: y = 16'hfe00;
			16'ha6e5: y = 16'hfe00;
			16'ha6e6: y = 16'hfe00;
			16'ha6e7: y = 16'hfe00;
			16'ha6e8: y = 16'hfe00;
			16'ha6e9: y = 16'hfe00;
			16'ha6ea: y = 16'hfe00;
			16'ha6eb: y = 16'hfe00;
			16'ha6ec: y = 16'hfe00;
			16'ha6ed: y = 16'hfe00;
			16'ha6ee: y = 16'hfe00;
			16'ha6ef: y = 16'hfe00;
			16'ha6f0: y = 16'hfe00;
			16'ha6f1: y = 16'hfe00;
			16'ha6f2: y = 16'hfe00;
			16'ha6f3: y = 16'hfe00;
			16'ha6f4: y = 16'hfe00;
			16'ha6f5: y = 16'hfe00;
			16'ha6f6: y = 16'hfe00;
			16'ha6f7: y = 16'hfe00;
			16'ha6f8: y = 16'hfe00;
			16'ha6f9: y = 16'hfe00;
			16'ha6fa: y = 16'hfe00;
			16'ha6fb: y = 16'hfe00;
			16'ha6fc: y = 16'hfe00;
			16'ha6fd: y = 16'hfe00;
			16'ha6fe: y = 16'hfe00;
			16'ha6ff: y = 16'hfe00;
			16'ha700: y = 16'hfe00;
			16'ha701: y = 16'hfe00;
			16'ha702: y = 16'hfe00;
			16'ha703: y = 16'hfe00;
			16'ha704: y = 16'hfe00;
			16'ha705: y = 16'hfe00;
			16'ha706: y = 16'hfe00;
			16'ha707: y = 16'hfe00;
			16'ha708: y = 16'hfe00;
			16'ha709: y = 16'hfe00;
			16'ha70a: y = 16'hfe00;
			16'ha70b: y = 16'hfe00;
			16'ha70c: y = 16'hfe00;
			16'ha70d: y = 16'hfe00;
			16'ha70e: y = 16'hfe00;
			16'ha70f: y = 16'hfe00;
			16'ha710: y = 16'hfe00;
			16'ha711: y = 16'hfe00;
			16'ha712: y = 16'hfe00;
			16'ha713: y = 16'hfe00;
			16'ha714: y = 16'hfe00;
			16'ha715: y = 16'hfe00;
			16'ha716: y = 16'hfe00;
			16'ha717: y = 16'hfe00;
			16'ha718: y = 16'hfe00;
			16'ha719: y = 16'hfe00;
			16'ha71a: y = 16'hfe00;
			16'ha71b: y = 16'hfe00;
			16'ha71c: y = 16'hfe00;
			16'ha71d: y = 16'hfe00;
			16'ha71e: y = 16'hfe00;
			16'ha71f: y = 16'hfe00;
			16'ha720: y = 16'hfe00;
			16'ha721: y = 16'hfe00;
			16'ha722: y = 16'hfe00;
			16'ha723: y = 16'hfe00;
			16'ha724: y = 16'hfe00;
			16'ha725: y = 16'hfe00;
			16'ha726: y = 16'hfe00;
			16'ha727: y = 16'hfe00;
			16'ha728: y = 16'hfe00;
			16'ha729: y = 16'hfe00;
			16'ha72a: y = 16'hfe00;
			16'ha72b: y = 16'hfe00;
			16'ha72c: y = 16'hfe00;
			16'ha72d: y = 16'hfe00;
			16'ha72e: y = 16'hfe00;
			16'ha72f: y = 16'hfe00;
			16'ha730: y = 16'hfe00;
			16'ha731: y = 16'hfe00;
			16'ha732: y = 16'hfe00;
			16'ha733: y = 16'hfe00;
			16'ha734: y = 16'hfe00;
			16'ha735: y = 16'hfe00;
			16'ha736: y = 16'hfe00;
			16'ha737: y = 16'hfe00;
			16'ha738: y = 16'hfe00;
			16'ha739: y = 16'hfe00;
			16'ha73a: y = 16'hfe00;
			16'ha73b: y = 16'hfe00;
			16'ha73c: y = 16'hfe00;
			16'ha73d: y = 16'hfe00;
			16'ha73e: y = 16'hfe00;
			16'ha73f: y = 16'hfe00;
			16'ha740: y = 16'hfe00;
			16'ha741: y = 16'hfe00;
			16'ha742: y = 16'hfe00;
			16'ha743: y = 16'hfe00;
			16'ha744: y = 16'hfe00;
			16'ha745: y = 16'hfe00;
			16'ha746: y = 16'hfe00;
			16'ha747: y = 16'hfe00;
			16'ha748: y = 16'hfe00;
			16'ha749: y = 16'hfe00;
			16'ha74a: y = 16'hfe00;
			16'ha74b: y = 16'hfe00;
			16'ha74c: y = 16'hfe00;
			16'ha74d: y = 16'hfe00;
			16'ha74e: y = 16'hfe00;
			16'ha74f: y = 16'hfe00;
			16'ha750: y = 16'hfe00;
			16'ha751: y = 16'hfe00;
			16'ha752: y = 16'hfe00;
			16'ha753: y = 16'hfe00;
			16'ha754: y = 16'hfe00;
			16'ha755: y = 16'hfe00;
			16'ha756: y = 16'hfe00;
			16'ha757: y = 16'hfe00;
			16'ha758: y = 16'hfe00;
			16'ha759: y = 16'hfe00;
			16'ha75a: y = 16'hfe00;
			16'ha75b: y = 16'hfe00;
			16'ha75c: y = 16'hfe00;
			16'ha75d: y = 16'hfe00;
			16'ha75e: y = 16'hfe00;
			16'ha75f: y = 16'hfe00;
			16'ha760: y = 16'hfe00;
			16'ha761: y = 16'hfe00;
			16'ha762: y = 16'hfe00;
			16'ha763: y = 16'hfe00;
			16'ha764: y = 16'hfe00;
			16'ha765: y = 16'hfe00;
			16'ha766: y = 16'hfe00;
			16'ha767: y = 16'hfe00;
			16'ha768: y = 16'hfe00;
			16'ha769: y = 16'hfe00;
			16'ha76a: y = 16'hfe00;
			16'ha76b: y = 16'hfe00;
			16'ha76c: y = 16'hfe00;
			16'ha76d: y = 16'hfe00;
			16'ha76e: y = 16'hfe00;
			16'ha76f: y = 16'hfe00;
			16'ha770: y = 16'hfe00;
			16'ha771: y = 16'hfe00;
			16'ha772: y = 16'hfe00;
			16'ha773: y = 16'hfe00;
			16'ha774: y = 16'hfe00;
			16'ha775: y = 16'hfe00;
			16'ha776: y = 16'hfe00;
			16'ha777: y = 16'hfe00;
			16'ha778: y = 16'hfe00;
			16'ha779: y = 16'hfe00;
			16'ha77a: y = 16'hfe00;
			16'ha77b: y = 16'hfe00;
			16'ha77c: y = 16'hfe00;
			16'ha77d: y = 16'hfe00;
			16'ha77e: y = 16'hfe00;
			16'ha77f: y = 16'hfe00;
			16'ha780: y = 16'hfe00;
			16'ha781: y = 16'hfe00;
			16'ha782: y = 16'hfe00;
			16'ha783: y = 16'hfe00;
			16'ha784: y = 16'hfe00;
			16'ha785: y = 16'hfe00;
			16'ha786: y = 16'hfe00;
			16'ha787: y = 16'hfe00;
			16'ha788: y = 16'hfe00;
			16'ha789: y = 16'hfe00;
			16'ha78a: y = 16'hfe00;
			16'ha78b: y = 16'hfe00;
			16'ha78c: y = 16'hfe00;
			16'ha78d: y = 16'hfe00;
			16'ha78e: y = 16'hfe00;
			16'ha78f: y = 16'hfe00;
			16'ha790: y = 16'hfe00;
			16'ha791: y = 16'hfe00;
			16'ha792: y = 16'hfe00;
			16'ha793: y = 16'hfe00;
			16'ha794: y = 16'hfe00;
			16'ha795: y = 16'hfe00;
			16'ha796: y = 16'hfe00;
			16'ha797: y = 16'hfe00;
			16'ha798: y = 16'hfe00;
			16'ha799: y = 16'hfe00;
			16'ha79a: y = 16'hfe00;
			16'ha79b: y = 16'hfe00;
			16'ha79c: y = 16'hfe00;
			16'ha79d: y = 16'hfe00;
			16'ha79e: y = 16'hfe00;
			16'ha79f: y = 16'hfe00;
			16'ha7a0: y = 16'hfe00;
			16'ha7a1: y = 16'hfe00;
			16'ha7a2: y = 16'hfe00;
			16'ha7a3: y = 16'hfe00;
			16'ha7a4: y = 16'hfe00;
			16'ha7a5: y = 16'hfe00;
			16'ha7a6: y = 16'hfe00;
			16'ha7a7: y = 16'hfe00;
			16'ha7a8: y = 16'hfe00;
			16'ha7a9: y = 16'hfe00;
			16'ha7aa: y = 16'hfe00;
			16'ha7ab: y = 16'hfe00;
			16'ha7ac: y = 16'hfe00;
			16'ha7ad: y = 16'hfe00;
			16'ha7ae: y = 16'hfe00;
			16'ha7af: y = 16'hfe00;
			16'ha7b0: y = 16'hfe00;
			16'ha7b1: y = 16'hfe00;
			16'ha7b2: y = 16'hfe00;
			16'ha7b3: y = 16'hfe00;
			16'ha7b4: y = 16'hfe00;
			16'ha7b5: y = 16'hfe00;
			16'ha7b6: y = 16'hfe00;
			16'ha7b7: y = 16'hfe00;
			16'ha7b8: y = 16'hfe00;
			16'ha7b9: y = 16'hfe00;
			16'ha7ba: y = 16'hfe00;
			16'ha7bb: y = 16'hfe00;
			16'ha7bc: y = 16'hfe00;
			16'ha7bd: y = 16'hfe00;
			16'ha7be: y = 16'hfe00;
			16'ha7bf: y = 16'hfe00;
			16'ha7c0: y = 16'hfe00;
			16'ha7c1: y = 16'hfe00;
			16'ha7c2: y = 16'hfe00;
			16'ha7c3: y = 16'hfe00;
			16'ha7c4: y = 16'hfe00;
			16'ha7c5: y = 16'hfe00;
			16'ha7c6: y = 16'hfe00;
			16'ha7c7: y = 16'hfe00;
			16'ha7c8: y = 16'hfe00;
			16'ha7c9: y = 16'hfe00;
			16'ha7ca: y = 16'hfe00;
			16'ha7cb: y = 16'hfe00;
			16'ha7cc: y = 16'hfe00;
			16'ha7cd: y = 16'hfe00;
			16'ha7ce: y = 16'hfe00;
			16'ha7cf: y = 16'hfe00;
			16'ha7d0: y = 16'hfe00;
			16'ha7d1: y = 16'hfe00;
			16'ha7d2: y = 16'hfe00;
			16'ha7d3: y = 16'hfe00;
			16'ha7d4: y = 16'hfe00;
			16'ha7d5: y = 16'hfe00;
			16'ha7d6: y = 16'hfe00;
			16'ha7d7: y = 16'hfe00;
			16'ha7d8: y = 16'hfe00;
			16'ha7d9: y = 16'hfe00;
			16'ha7da: y = 16'hfe00;
			16'ha7db: y = 16'hfe00;
			16'ha7dc: y = 16'hfe00;
			16'ha7dd: y = 16'hfe00;
			16'ha7de: y = 16'hfe00;
			16'ha7df: y = 16'hfe00;
			16'ha7e0: y = 16'hfe00;
			16'ha7e1: y = 16'hfe00;
			16'ha7e2: y = 16'hfe00;
			16'ha7e3: y = 16'hfe00;
			16'ha7e4: y = 16'hfe00;
			16'ha7e5: y = 16'hfe00;
			16'ha7e6: y = 16'hfe00;
			16'ha7e7: y = 16'hfe00;
			16'ha7e8: y = 16'hfe00;
			16'ha7e9: y = 16'hfe00;
			16'ha7ea: y = 16'hfe00;
			16'ha7eb: y = 16'hfe00;
			16'ha7ec: y = 16'hfe00;
			16'ha7ed: y = 16'hfe00;
			16'ha7ee: y = 16'hfe00;
			16'ha7ef: y = 16'hfe00;
			16'ha7f0: y = 16'hfe00;
			16'ha7f1: y = 16'hfe00;
			16'ha7f2: y = 16'hfe00;
			16'ha7f3: y = 16'hfe00;
			16'ha7f4: y = 16'hfe00;
			16'ha7f5: y = 16'hfe00;
			16'ha7f6: y = 16'hfe00;
			16'ha7f7: y = 16'hfe00;
			16'ha7f8: y = 16'hfe00;
			16'ha7f9: y = 16'hfe00;
			16'ha7fa: y = 16'hfe00;
			16'ha7fb: y = 16'hfe00;
			16'ha7fc: y = 16'hfe00;
			16'ha7fd: y = 16'hfe00;
			16'ha7fe: y = 16'hfe00;
			16'ha7ff: y = 16'hfe00;
			16'ha800: y = 16'hfe00;
			16'ha801: y = 16'hfe00;
			16'ha802: y = 16'hfe00;
			16'ha803: y = 16'hfe00;
			16'ha804: y = 16'hfe00;
			16'ha805: y = 16'hfe00;
			16'ha806: y = 16'hfe00;
			16'ha807: y = 16'hfe00;
			16'ha808: y = 16'hfe00;
			16'ha809: y = 16'hfe00;
			16'ha80a: y = 16'hfe00;
			16'ha80b: y = 16'hfe00;
			16'ha80c: y = 16'hfe00;
			16'ha80d: y = 16'hfe00;
			16'ha80e: y = 16'hfe00;
			16'ha80f: y = 16'hfe00;
			16'ha810: y = 16'hfe00;
			16'ha811: y = 16'hfe00;
			16'ha812: y = 16'hfe00;
			16'ha813: y = 16'hfe00;
			16'ha814: y = 16'hfe00;
			16'ha815: y = 16'hfe00;
			16'ha816: y = 16'hfe00;
			16'ha817: y = 16'hfe00;
			16'ha818: y = 16'hfe00;
			16'ha819: y = 16'hfe00;
			16'ha81a: y = 16'hfe00;
			16'ha81b: y = 16'hfe00;
			16'ha81c: y = 16'hfe00;
			16'ha81d: y = 16'hfe00;
			16'ha81e: y = 16'hfe00;
			16'ha81f: y = 16'hfe00;
			16'ha820: y = 16'hfe00;
			16'ha821: y = 16'hfe00;
			16'ha822: y = 16'hfe00;
			16'ha823: y = 16'hfe00;
			16'ha824: y = 16'hfe00;
			16'ha825: y = 16'hfe00;
			16'ha826: y = 16'hfe00;
			16'ha827: y = 16'hfe00;
			16'ha828: y = 16'hfe00;
			16'ha829: y = 16'hfe00;
			16'ha82a: y = 16'hfe00;
			16'ha82b: y = 16'hfe00;
			16'ha82c: y = 16'hfe00;
			16'ha82d: y = 16'hfe00;
			16'ha82e: y = 16'hfe00;
			16'ha82f: y = 16'hfe00;
			16'ha830: y = 16'hfe00;
			16'ha831: y = 16'hfe00;
			16'ha832: y = 16'hfe00;
			16'ha833: y = 16'hfe00;
			16'ha834: y = 16'hfe00;
			16'ha835: y = 16'hfe00;
			16'ha836: y = 16'hfe00;
			16'ha837: y = 16'hfe00;
			16'ha838: y = 16'hfe00;
			16'ha839: y = 16'hfe00;
			16'ha83a: y = 16'hfe00;
			16'ha83b: y = 16'hfe00;
			16'ha83c: y = 16'hfe00;
			16'ha83d: y = 16'hfe00;
			16'ha83e: y = 16'hfe00;
			16'ha83f: y = 16'hfe00;
			16'ha840: y = 16'hfe00;
			16'ha841: y = 16'hfe00;
			16'ha842: y = 16'hfe00;
			16'ha843: y = 16'hfe00;
			16'ha844: y = 16'hfe00;
			16'ha845: y = 16'hfe00;
			16'ha846: y = 16'hfe00;
			16'ha847: y = 16'hfe00;
			16'ha848: y = 16'hfe00;
			16'ha849: y = 16'hfe00;
			16'ha84a: y = 16'hfe00;
			16'ha84b: y = 16'hfe00;
			16'ha84c: y = 16'hfe00;
			16'ha84d: y = 16'hfe00;
			16'ha84e: y = 16'hfe00;
			16'ha84f: y = 16'hfe00;
			16'ha850: y = 16'hfe00;
			16'ha851: y = 16'hfe00;
			16'ha852: y = 16'hfe00;
			16'ha853: y = 16'hfe00;
			16'ha854: y = 16'hfe00;
			16'ha855: y = 16'hfe00;
			16'ha856: y = 16'hfe00;
			16'ha857: y = 16'hfe00;
			16'ha858: y = 16'hfe00;
			16'ha859: y = 16'hfe00;
			16'ha85a: y = 16'hfe00;
			16'ha85b: y = 16'hfe00;
			16'ha85c: y = 16'hfe00;
			16'ha85d: y = 16'hfe00;
			16'ha85e: y = 16'hfe00;
			16'ha85f: y = 16'hfe00;
			16'ha860: y = 16'hfe00;
			16'ha861: y = 16'hfe00;
			16'ha862: y = 16'hfe00;
			16'ha863: y = 16'hfe00;
			16'ha864: y = 16'hfe00;
			16'ha865: y = 16'hfe00;
			16'ha866: y = 16'hfe00;
			16'ha867: y = 16'hfe00;
			16'ha868: y = 16'hfe00;
			16'ha869: y = 16'hfe00;
			16'ha86a: y = 16'hfe00;
			16'ha86b: y = 16'hfe00;
			16'ha86c: y = 16'hfe00;
			16'ha86d: y = 16'hfe00;
			16'ha86e: y = 16'hfe00;
			16'ha86f: y = 16'hfe00;
			16'ha870: y = 16'hfe00;
			16'ha871: y = 16'hfe00;
			16'ha872: y = 16'hfe00;
			16'ha873: y = 16'hfe00;
			16'ha874: y = 16'hfe00;
			16'ha875: y = 16'hfe00;
			16'ha876: y = 16'hfe00;
			16'ha877: y = 16'hfe00;
			16'ha878: y = 16'hfe00;
			16'ha879: y = 16'hfe00;
			16'ha87a: y = 16'hfe00;
			16'ha87b: y = 16'hfe00;
			16'ha87c: y = 16'hfe00;
			16'ha87d: y = 16'hfe00;
			16'ha87e: y = 16'hfe00;
			16'ha87f: y = 16'hfe00;
			16'ha880: y = 16'hfe00;
			16'ha881: y = 16'hfe00;
			16'ha882: y = 16'hfe00;
			16'ha883: y = 16'hfe00;
			16'ha884: y = 16'hfe00;
			16'ha885: y = 16'hfe00;
			16'ha886: y = 16'hfe00;
			16'ha887: y = 16'hfe00;
			16'ha888: y = 16'hfe00;
			16'ha889: y = 16'hfe00;
			16'ha88a: y = 16'hfe00;
			16'ha88b: y = 16'hfe00;
			16'ha88c: y = 16'hfe00;
			16'ha88d: y = 16'hfe00;
			16'ha88e: y = 16'hfe00;
			16'ha88f: y = 16'hfe00;
			16'ha890: y = 16'hfe00;
			16'ha891: y = 16'hfe00;
			16'ha892: y = 16'hfe00;
			16'ha893: y = 16'hfe00;
			16'ha894: y = 16'hfe00;
			16'ha895: y = 16'hfe00;
			16'ha896: y = 16'hfe00;
			16'ha897: y = 16'hfe00;
			16'ha898: y = 16'hfe00;
			16'ha899: y = 16'hfe00;
			16'ha89a: y = 16'hfe00;
			16'ha89b: y = 16'hfe00;
			16'ha89c: y = 16'hfe00;
			16'ha89d: y = 16'hfe00;
			16'ha89e: y = 16'hfe00;
			16'ha89f: y = 16'hfe00;
			16'ha8a0: y = 16'hfe00;
			16'ha8a1: y = 16'hfe00;
			16'ha8a2: y = 16'hfe00;
			16'ha8a3: y = 16'hfe00;
			16'ha8a4: y = 16'hfe00;
			16'ha8a5: y = 16'hfe00;
			16'ha8a6: y = 16'hfe00;
			16'ha8a7: y = 16'hfe00;
			16'ha8a8: y = 16'hfe00;
			16'ha8a9: y = 16'hfe00;
			16'ha8aa: y = 16'hfe00;
			16'ha8ab: y = 16'hfe00;
			16'ha8ac: y = 16'hfe00;
			16'ha8ad: y = 16'hfe00;
			16'ha8ae: y = 16'hfe00;
			16'ha8af: y = 16'hfe00;
			16'ha8b0: y = 16'hfe00;
			16'ha8b1: y = 16'hfe00;
			16'ha8b2: y = 16'hfe00;
			16'ha8b3: y = 16'hfe00;
			16'ha8b4: y = 16'hfe00;
			16'ha8b5: y = 16'hfe00;
			16'ha8b6: y = 16'hfe00;
			16'ha8b7: y = 16'hfe00;
			16'ha8b8: y = 16'hfe00;
			16'ha8b9: y = 16'hfe00;
			16'ha8ba: y = 16'hfe00;
			16'ha8bb: y = 16'hfe00;
			16'ha8bc: y = 16'hfe00;
			16'ha8bd: y = 16'hfe00;
			16'ha8be: y = 16'hfe00;
			16'ha8bf: y = 16'hfe00;
			16'ha8c0: y = 16'hfe00;
			16'ha8c1: y = 16'hfe00;
			16'ha8c2: y = 16'hfe00;
			16'ha8c3: y = 16'hfe00;
			16'ha8c4: y = 16'hfe00;
			16'ha8c5: y = 16'hfe00;
			16'ha8c6: y = 16'hfe00;
			16'ha8c7: y = 16'hfe00;
			16'ha8c8: y = 16'hfe00;
			16'ha8c9: y = 16'hfe00;
			16'ha8ca: y = 16'hfe00;
			16'ha8cb: y = 16'hfe00;
			16'ha8cc: y = 16'hfe00;
			16'ha8cd: y = 16'hfe00;
			16'ha8ce: y = 16'hfe00;
			16'ha8cf: y = 16'hfe00;
			16'ha8d0: y = 16'hfe00;
			16'ha8d1: y = 16'hfe00;
			16'ha8d2: y = 16'hfe00;
			16'ha8d3: y = 16'hfe00;
			16'ha8d4: y = 16'hfe00;
			16'ha8d5: y = 16'hfe00;
			16'ha8d6: y = 16'hfe00;
			16'ha8d7: y = 16'hfe00;
			16'ha8d8: y = 16'hfe00;
			16'ha8d9: y = 16'hfe00;
			16'ha8da: y = 16'hfe00;
			16'ha8db: y = 16'hfe00;
			16'ha8dc: y = 16'hfe00;
			16'ha8dd: y = 16'hfe00;
			16'ha8de: y = 16'hfe00;
			16'ha8df: y = 16'hfe00;
			16'ha8e0: y = 16'hfe00;
			16'ha8e1: y = 16'hfe00;
			16'ha8e2: y = 16'hfe00;
			16'ha8e3: y = 16'hfe00;
			16'ha8e4: y = 16'hfe00;
			16'ha8e5: y = 16'hfe00;
			16'ha8e6: y = 16'hfe00;
			16'ha8e7: y = 16'hfe00;
			16'ha8e8: y = 16'hfe00;
			16'ha8e9: y = 16'hfe00;
			16'ha8ea: y = 16'hfe00;
			16'ha8eb: y = 16'hfe00;
			16'ha8ec: y = 16'hfe00;
			16'ha8ed: y = 16'hfe00;
			16'ha8ee: y = 16'hfe00;
			16'ha8ef: y = 16'hfe00;
			16'ha8f0: y = 16'hfe00;
			16'ha8f1: y = 16'hfe00;
			16'ha8f2: y = 16'hfe00;
			16'ha8f3: y = 16'hfe00;
			16'ha8f4: y = 16'hfe00;
			16'ha8f5: y = 16'hfe00;
			16'ha8f6: y = 16'hfe00;
			16'ha8f7: y = 16'hfe00;
			16'ha8f8: y = 16'hfe00;
			16'ha8f9: y = 16'hfe00;
			16'ha8fa: y = 16'hfe00;
			16'ha8fb: y = 16'hfe00;
			16'ha8fc: y = 16'hfe00;
			16'ha8fd: y = 16'hfe00;
			16'ha8fe: y = 16'hfe00;
			16'ha8ff: y = 16'hfe00;
			16'ha900: y = 16'hfe00;
			16'ha901: y = 16'hfe00;
			16'ha902: y = 16'hfe00;
			16'ha903: y = 16'hfe00;
			16'ha904: y = 16'hfe00;
			16'ha905: y = 16'hfe00;
			16'ha906: y = 16'hfe00;
			16'ha907: y = 16'hfe00;
			16'ha908: y = 16'hfe00;
			16'ha909: y = 16'hfe00;
			16'ha90a: y = 16'hfe00;
			16'ha90b: y = 16'hfe00;
			16'ha90c: y = 16'hfe00;
			16'ha90d: y = 16'hfe00;
			16'ha90e: y = 16'hfe00;
			16'ha90f: y = 16'hfe00;
			16'ha910: y = 16'hfe00;
			16'ha911: y = 16'hfe00;
			16'ha912: y = 16'hfe00;
			16'ha913: y = 16'hfe00;
			16'ha914: y = 16'hfe00;
			16'ha915: y = 16'hfe00;
			16'ha916: y = 16'hfe00;
			16'ha917: y = 16'hfe00;
			16'ha918: y = 16'hfe00;
			16'ha919: y = 16'hfe00;
			16'ha91a: y = 16'hfe00;
			16'ha91b: y = 16'hfe00;
			16'ha91c: y = 16'hfe00;
			16'ha91d: y = 16'hfe00;
			16'ha91e: y = 16'hfe00;
			16'ha91f: y = 16'hfe00;
			16'ha920: y = 16'hfe00;
			16'ha921: y = 16'hfe00;
			16'ha922: y = 16'hfe00;
			16'ha923: y = 16'hfe00;
			16'ha924: y = 16'hfe00;
			16'ha925: y = 16'hfe00;
			16'ha926: y = 16'hfe00;
			16'ha927: y = 16'hfe00;
			16'ha928: y = 16'hfe00;
			16'ha929: y = 16'hfe00;
			16'ha92a: y = 16'hfe00;
			16'ha92b: y = 16'hfe00;
			16'ha92c: y = 16'hfe00;
			16'ha92d: y = 16'hfe00;
			16'ha92e: y = 16'hfe00;
			16'ha92f: y = 16'hfe00;
			16'ha930: y = 16'hfe00;
			16'ha931: y = 16'hfe00;
			16'ha932: y = 16'hfe00;
			16'ha933: y = 16'hfe00;
			16'ha934: y = 16'hfe00;
			16'ha935: y = 16'hfe00;
			16'ha936: y = 16'hfe00;
			16'ha937: y = 16'hfe00;
			16'ha938: y = 16'hfe00;
			16'ha939: y = 16'hfe00;
			16'ha93a: y = 16'hfe00;
			16'ha93b: y = 16'hfe00;
			16'ha93c: y = 16'hfe00;
			16'ha93d: y = 16'hfe00;
			16'ha93e: y = 16'hfe00;
			16'ha93f: y = 16'hfe00;
			16'ha940: y = 16'hfe00;
			16'ha941: y = 16'hfe00;
			16'ha942: y = 16'hfe00;
			16'ha943: y = 16'hfe00;
			16'ha944: y = 16'hfe00;
			16'ha945: y = 16'hfe00;
			16'ha946: y = 16'hfe00;
			16'ha947: y = 16'hfe00;
			16'ha948: y = 16'hfe00;
			16'ha949: y = 16'hfe00;
			16'ha94a: y = 16'hfe00;
			16'ha94b: y = 16'hfe00;
			16'ha94c: y = 16'hfe00;
			16'ha94d: y = 16'hfe00;
			16'ha94e: y = 16'hfe00;
			16'ha94f: y = 16'hfe00;
			16'ha950: y = 16'hfe00;
			16'ha951: y = 16'hfe00;
			16'ha952: y = 16'hfe00;
			16'ha953: y = 16'hfe00;
			16'ha954: y = 16'hfe00;
			16'ha955: y = 16'hfe00;
			16'ha956: y = 16'hfe00;
			16'ha957: y = 16'hfe00;
			16'ha958: y = 16'hfe00;
			16'ha959: y = 16'hfe00;
			16'ha95a: y = 16'hfe00;
			16'ha95b: y = 16'hfe00;
			16'ha95c: y = 16'hfe00;
			16'ha95d: y = 16'hfe00;
			16'ha95e: y = 16'hfe00;
			16'ha95f: y = 16'hfe00;
			16'ha960: y = 16'hfe00;
			16'ha961: y = 16'hfe00;
			16'ha962: y = 16'hfe00;
			16'ha963: y = 16'hfe00;
			16'ha964: y = 16'hfe00;
			16'ha965: y = 16'hfe00;
			16'ha966: y = 16'hfe00;
			16'ha967: y = 16'hfe00;
			16'ha968: y = 16'hfe00;
			16'ha969: y = 16'hfe00;
			16'ha96a: y = 16'hfe00;
			16'ha96b: y = 16'hfe00;
			16'ha96c: y = 16'hfe00;
			16'ha96d: y = 16'hfe00;
			16'ha96e: y = 16'hfe00;
			16'ha96f: y = 16'hfe00;
			16'ha970: y = 16'hfe00;
			16'ha971: y = 16'hfe00;
			16'ha972: y = 16'hfe00;
			16'ha973: y = 16'hfe00;
			16'ha974: y = 16'hfe00;
			16'ha975: y = 16'hfe00;
			16'ha976: y = 16'hfe00;
			16'ha977: y = 16'hfe00;
			16'ha978: y = 16'hfe00;
			16'ha979: y = 16'hfe00;
			16'ha97a: y = 16'hfe00;
			16'ha97b: y = 16'hfe00;
			16'ha97c: y = 16'hfe00;
			16'ha97d: y = 16'hfe00;
			16'ha97e: y = 16'hfe00;
			16'ha97f: y = 16'hfe00;
			16'ha980: y = 16'hfe00;
			16'ha981: y = 16'hfe00;
			16'ha982: y = 16'hfe00;
			16'ha983: y = 16'hfe00;
			16'ha984: y = 16'hfe00;
			16'ha985: y = 16'hfe00;
			16'ha986: y = 16'hfe00;
			16'ha987: y = 16'hfe00;
			16'ha988: y = 16'hfe00;
			16'ha989: y = 16'hfe00;
			16'ha98a: y = 16'hfe00;
			16'ha98b: y = 16'hfe00;
			16'ha98c: y = 16'hfe00;
			16'ha98d: y = 16'hfe00;
			16'ha98e: y = 16'hfe00;
			16'ha98f: y = 16'hfe00;
			16'ha990: y = 16'hfe00;
			16'ha991: y = 16'hfe00;
			16'ha992: y = 16'hfe00;
			16'ha993: y = 16'hfe00;
			16'ha994: y = 16'hfe00;
			16'ha995: y = 16'hfe00;
			16'ha996: y = 16'hfe00;
			16'ha997: y = 16'hfe00;
			16'ha998: y = 16'hfe00;
			16'ha999: y = 16'hfe00;
			16'ha99a: y = 16'hfe00;
			16'ha99b: y = 16'hfe00;
			16'ha99c: y = 16'hfe00;
			16'ha99d: y = 16'hfe00;
			16'ha99e: y = 16'hfe00;
			16'ha99f: y = 16'hfe00;
			16'ha9a0: y = 16'hfe00;
			16'ha9a1: y = 16'hfe00;
			16'ha9a2: y = 16'hfe00;
			16'ha9a3: y = 16'hfe00;
			16'ha9a4: y = 16'hfe00;
			16'ha9a5: y = 16'hfe00;
			16'ha9a6: y = 16'hfe00;
			16'ha9a7: y = 16'hfe00;
			16'ha9a8: y = 16'hfe00;
			16'ha9a9: y = 16'hfe00;
			16'ha9aa: y = 16'hfe00;
			16'ha9ab: y = 16'hfe00;
			16'ha9ac: y = 16'hfe00;
			16'ha9ad: y = 16'hfe00;
			16'ha9ae: y = 16'hfe00;
			16'ha9af: y = 16'hfe00;
			16'ha9b0: y = 16'hfe00;
			16'ha9b1: y = 16'hfe00;
			16'ha9b2: y = 16'hfe00;
			16'ha9b3: y = 16'hfe00;
			16'ha9b4: y = 16'hfe00;
			16'ha9b5: y = 16'hfe00;
			16'ha9b6: y = 16'hfe00;
			16'ha9b7: y = 16'hfe00;
			16'ha9b8: y = 16'hfe00;
			16'ha9b9: y = 16'hfe00;
			16'ha9ba: y = 16'hfe00;
			16'ha9bb: y = 16'hfe00;
			16'ha9bc: y = 16'hfe00;
			16'ha9bd: y = 16'hfe00;
			16'ha9be: y = 16'hfe00;
			16'ha9bf: y = 16'hfe00;
			16'ha9c0: y = 16'hfe00;
			16'ha9c1: y = 16'hfe00;
			16'ha9c2: y = 16'hfe00;
			16'ha9c3: y = 16'hfe00;
			16'ha9c4: y = 16'hfe00;
			16'ha9c5: y = 16'hfe00;
			16'ha9c6: y = 16'hfe00;
			16'ha9c7: y = 16'hfe00;
			16'ha9c8: y = 16'hfe00;
			16'ha9c9: y = 16'hfe00;
			16'ha9ca: y = 16'hfe00;
			16'ha9cb: y = 16'hfe00;
			16'ha9cc: y = 16'hfe00;
			16'ha9cd: y = 16'hfe00;
			16'ha9ce: y = 16'hfe00;
			16'ha9cf: y = 16'hfe00;
			16'ha9d0: y = 16'hfe00;
			16'ha9d1: y = 16'hfe00;
			16'ha9d2: y = 16'hfe00;
			16'ha9d3: y = 16'hfe00;
			16'ha9d4: y = 16'hfe00;
			16'ha9d5: y = 16'hfe00;
			16'ha9d6: y = 16'hfe00;
			16'ha9d7: y = 16'hfe00;
			16'ha9d8: y = 16'hfe00;
			16'ha9d9: y = 16'hfe00;
			16'ha9da: y = 16'hfe00;
			16'ha9db: y = 16'hfe00;
			16'ha9dc: y = 16'hfe00;
			16'ha9dd: y = 16'hfe00;
			16'ha9de: y = 16'hfe00;
			16'ha9df: y = 16'hfe00;
			16'ha9e0: y = 16'hfe00;
			16'ha9e1: y = 16'hfe00;
			16'ha9e2: y = 16'hfe00;
			16'ha9e3: y = 16'hfe00;
			16'ha9e4: y = 16'hfe00;
			16'ha9e5: y = 16'hfe00;
			16'ha9e6: y = 16'hfe00;
			16'ha9e7: y = 16'hfe00;
			16'ha9e8: y = 16'hfe00;
			16'ha9e9: y = 16'hfe00;
			16'ha9ea: y = 16'hfe00;
			16'ha9eb: y = 16'hfe00;
			16'ha9ec: y = 16'hfe00;
			16'ha9ed: y = 16'hfe00;
			16'ha9ee: y = 16'hfe00;
			16'ha9ef: y = 16'hfe00;
			16'ha9f0: y = 16'hfe00;
			16'ha9f1: y = 16'hfe00;
			16'ha9f2: y = 16'hfe00;
			16'ha9f3: y = 16'hfe00;
			16'ha9f4: y = 16'hfe00;
			16'ha9f5: y = 16'hfe00;
			16'ha9f6: y = 16'hfe00;
			16'ha9f7: y = 16'hfe00;
			16'ha9f8: y = 16'hfe00;
			16'ha9f9: y = 16'hfe00;
			16'ha9fa: y = 16'hfe00;
			16'ha9fb: y = 16'hfe00;
			16'ha9fc: y = 16'hfe00;
			16'ha9fd: y = 16'hfe00;
			16'ha9fe: y = 16'hfe00;
			16'ha9ff: y = 16'hfe00;
			16'haa00: y = 16'hfe00;
			16'haa01: y = 16'hfe00;
			16'haa02: y = 16'hfe00;
			16'haa03: y = 16'hfe00;
			16'haa04: y = 16'hfe00;
			16'haa05: y = 16'hfe00;
			16'haa06: y = 16'hfe00;
			16'haa07: y = 16'hfe00;
			16'haa08: y = 16'hfe00;
			16'haa09: y = 16'hfe00;
			16'haa0a: y = 16'hfe00;
			16'haa0b: y = 16'hfe00;
			16'haa0c: y = 16'hfe00;
			16'haa0d: y = 16'hfe00;
			16'haa0e: y = 16'hfe00;
			16'haa0f: y = 16'hfe00;
			16'haa10: y = 16'hfe00;
			16'haa11: y = 16'hfe00;
			16'haa12: y = 16'hfe00;
			16'haa13: y = 16'hfe00;
			16'haa14: y = 16'hfe00;
			16'haa15: y = 16'hfe00;
			16'haa16: y = 16'hfe00;
			16'haa17: y = 16'hfe00;
			16'haa18: y = 16'hfe00;
			16'haa19: y = 16'hfe00;
			16'haa1a: y = 16'hfe00;
			16'haa1b: y = 16'hfe00;
			16'haa1c: y = 16'hfe00;
			16'haa1d: y = 16'hfe00;
			16'haa1e: y = 16'hfe00;
			16'haa1f: y = 16'hfe00;
			16'haa20: y = 16'hfe00;
			16'haa21: y = 16'hfe00;
			16'haa22: y = 16'hfe00;
			16'haa23: y = 16'hfe00;
			16'haa24: y = 16'hfe00;
			16'haa25: y = 16'hfe00;
			16'haa26: y = 16'hfe00;
			16'haa27: y = 16'hfe00;
			16'haa28: y = 16'hfe00;
			16'haa29: y = 16'hfe00;
			16'haa2a: y = 16'hfe00;
			16'haa2b: y = 16'hfe00;
			16'haa2c: y = 16'hfe00;
			16'haa2d: y = 16'hfe00;
			16'haa2e: y = 16'hfe00;
			16'haa2f: y = 16'hfe00;
			16'haa30: y = 16'hfe00;
			16'haa31: y = 16'hfe00;
			16'haa32: y = 16'hfe00;
			16'haa33: y = 16'hfe00;
			16'haa34: y = 16'hfe00;
			16'haa35: y = 16'hfe00;
			16'haa36: y = 16'hfe00;
			16'haa37: y = 16'hfe00;
			16'haa38: y = 16'hfe00;
			16'haa39: y = 16'hfe00;
			16'haa3a: y = 16'hfe00;
			16'haa3b: y = 16'hfe00;
			16'haa3c: y = 16'hfe00;
			16'haa3d: y = 16'hfe00;
			16'haa3e: y = 16'hfe00;
			16'haa3f: y = 16'hfe00;
			16'haa40: y = 16'hfe00;
			16'haa41: y = 16'hfe00;
			16'haa42: y = 16'hfe00;
			16'haa43: y = 16'hfe00;
			16'haa44: y = 16'hfe00;
			16'haa45: y = 16'hfe00;
			16'haa46: y = 16'hfe00;
			16'haa47: y = 16'hfe00;
			16'haa48: y = 16'hfe00;
			16'haa49: y = 16'hfe00;
			16'haa4a: y = 16'hfe00;
			16'haa4b: y = 16'hfe00;
			16'haa4c: y = 16'hfe00;
			16'haa4d: y = 16'hfe00;
			16'haa4e: y = 16'hfe00;
			16'haa4f: y = 16'hfe00;
			16'haa50: y = 16'hfe00;
			16'haa51: y = 16'hfe00;
			16'haa52: y = 16'hfe00;
			16'haa53: y = 16'hfe00;
			16'haa54: y = 16'hfe00;
			16'haa55: y = 16'hfe00;
			16'haa56: y = 16'hfe00;
			16'haa57: y = 16'hfe00;
			16'haa58: y = 16'hfe00;
			16'haa59: y = 16'hfe00;
			16'haa5a: y = 16'hfe00;
			16'haa5b: y = 16'hfe00;
			16'haa5c: y = 16'hfe00;
			16'haa5d: y = 16'hfe00;
			16'haa5e: y = 16'hfe00;
			16'haa5f: y = 16'hfe00;
			16'haa60: y = 16'hfe00;
			16'haa61: y = 16'hfe00;
			16'haa62: y = 16'hfe00;
			16'haa63: y = 16'hfe00;
			16'haa64: y = 16'hfe00;
			16'haa65: y = 16'hfe00;
			16'haa66: y = 16'hfe00;
			16'haa67: y = 16'hfe00;
			16'haa68: y = 16'hfe00;
			16'haa69: y = 16'hfe00;
			16'haa6a: y = 16'hfe00;
			16'haa6b: y = 16'hfe00;
			16'haa6c: y = 16'hfe00;
			16'haa6d: y = 16'hfe00;
			16'haa6e: y = 16'hfe00;
			16'haa6f: y = 16'hfe00;
			16'haa70: y = 16'hfe00;
			16'haa71: y = 16'hfe00;
			16'haa72: y = 16'hfe00;
			16'haa73: y = 16'hfe00;
			16'haa74: y = 16'hfe00;
			16'haa75: y = 16'hfe00;
			16'haa76: y = 16'hfe00;
			16'haa77: y = 16'hfe00;
			16'haa78: y = 16'hfe00;
			16'haa79: y = 16'hfe00;
			16'haa7a: y = 16'hfe00;
			16'haa7b: y = 16'hfe00;
			16'haa7c: y = 16'hfe00;
			16'haa7d: y = 16'hfe00;
			16'haa7e: y = 16'hfe00;
			16'haa7f: y = 16'hfe00;
			16'haa80: y = 16'hfe00;
			16'haa81: y = 16'hfe00;
			16'haa82: y = 16'hfe00;
			16'haa83: y = 16'hfe00;
			16'haa84: y = 16'hfe00;
			16'haa85: y = 16'hfe00;
			16'haa86: y = 16'hfe00;
			16'haa87: y = 16'hfe00;
			16'haa88: y = 16'hfe00;
			16'haa89: y = 16'hfe00;
			16'haa8a: y = 16'hfe00;
			16'haa8b: y = 16'hfe00;
			16'haa8c: y = 16'hfe00;
			16'haa8d: y = 16'hfe00;
			16'haa8e: y = 16'hfe00;
			16'haa8f: y = 16'hfe00;
			16'haa90: y = 16'hfe00;
			16'haa91: y = 16'hfe00;
			16'haa92: y = 16'hfe00;
			16'haa93: y = 16'hfe00;
			16'haa94: y = 16'hfe00;
			16'haa95: y = 16'hfe00;
			16'haa96: y = 16'hfe00;
			16'haa97: y = 16'hfe00;
			16'haa98: y = 16'hfe00;
			16'haa99: y = 16'hfe00;
			16'haa9a: y = 16'hfe00;
			16'haa9b: y = 16'hfe00;
			16'haa9c: y = 16'hfe00;
			16'haa9d: y = 16'hfe00;
			16'haa9e: y = 16'hfe00;
			16'haa9f: y = 16'hfe00;
			16'haaa0: y = 16'hfe00;
			16'haaa1: y = 16'hfe00;
			16'haaa2: y = 16'hfe00;
			16'haaa3: y = 16'hfe00;
			16'haaa4: y = 16'hfe00;
			16'haaa5: y = 16'hfe00;
			16'haaa6: y = 16'hfe00;
			16'haaa7: y = 16'hfe00;
			16'haaa8: y = 16'hfe00;
			16'haaa9: y = 16'hfe00;
			16'haaaa: y = 16'hfe00;
			16'haaab: y = 16'hfe00;
			16'haaac: y = 16'hfe00;
			16'haaad: y = 16'hfe00;
			16'haaae: y = 16'hfe00;
			16'haaaf: y = 16'hfe00;
			16'haab0: y = 16'hfe00;
			16'haab1: y = 16'hfe00;
			16'haab2: y = 16'hfe00;
			16'haab3: y = 16'hfe00;
			16'haab4: y = 16'hfe00;
			16'haab5: y = 16'hfe00;
			16'haab6: y = 16'hfe00;
			16'haab7: y = 16'hfe00;
			16'haab8: y = 16'hfe00;
			16'haab9: y = 16'hfe00;
			16'haaba: y = 16'hfe00;
			16'haabb: y = 16'hfe00;
			16'haabc: y = 16'hfe00;
			16'haabd: y = 16'hfe00;
			16'haabe: y = 16'hfe00;
			16'haabf: y = 16'hfe00;
			16'haac0: y = 16'hfe00;
			16'haac1: y = 16'hfe00;
			16'haac2: y = 16'hfe00;
			16'haac3: y = 16'hfe00;
			16'haac4: y = 16'hfe00;
			16'haac5: y = 16'hfe00;
			16'haac6: y = 16'hfe00;
			16'haac7: y = 16'hfe00;
			16'haac8: y = 16'hfe00;
			16'haac9: y = 16'hfe00;
			16'haaca: y = 16'hfe00;
			16'haacb: y = 16'hfe00;
			16'haacc: y = 16'hfe00;
			16'haacd: y = 16'hfe00;
			16'haace: y = 16'hfe00;
			16'haacf: y = 16'hfe00;
			16'haad0: y = 16'hfe00;
			16'haad1: y = 16'hfe00;
			16'haad2: y = 16'hfe00;
			16'haad3: y = 16'hfe00;
			16'haad4: y = 16'hfe00;
			16'haad5: y = 16'hfe00;
			16'haad6: y = 16'hfe00;
			16'haad7: y = 16'hfe00;
			16'haad8: y = 16'hfe00;
			16'haad9: y = 16'hfe00;
			16'haada: y = 16'hfe00;
			16'haadb: y = 16'hfe00;
			16'haadc: y = 16'hfe00;
			16'haadd: y = 16'hfe00;
			16'haade: y = 16'hfe00;
			16'haadf: y = 16'hfe00;
			16'haae0: y = 16'hfe00;
			16'haae1: y = 16'hfe00;
			16'haae2: y = 16'hfe00;
			16'haae3: y = 16'hfe00;
			16'haae4: y = 16'hfe00;
			16'haae5: y = 16'hfe00;
			16'haae6: y = 16'hfe00;
			16'haae7: y = 16'hfe00;
			16'haae8: y = 16'hfe00;
			16'haae9: y = 16'hfe00;
			16'haaea: y = 16'hfe00;
			16'haaeb: y = 16'hfe00;
			16'haaec: y = 16'hfe00;
			16'haaed: y = 16'hfe00;
			16'haaee: y = 16'hfe00;
			16'haaef: y = 16'hfe00;
			16'haaf0: y = 16'hfe00;
			16'haaf1: y = 16'hfe00;
			16'haaf2: y = 16'hfe00;
			16'haaf3: y = 16'hfe00;
			16'haaf4: y = 16'hfe00;
			16'haaf5: y = 16'hfe00;
			16'haaf6: y = 16'hfe00;
			16'haaf7: y = 16'hfe00;
			16'haaf8: y = 16'hfe00;
			16'haaf9: y = 16'hfe00;
			16'haafa: y = 16'hfe00;
			16'haafb: y = 16'hfe00;
			16'haafc: y = 16'hfe00;
			16'haafd: y = 16'hfe00;
			16'haafe: y = 16'hfe00;
			16'haaff: y = 16'hfe00;
			16'hab00: y = 16'hfe00;
			16'hab01: y = 16'hfe00;
			16'hab02: y = 16'hfe00;
			16'hab03: y = 16'hfe00;
			16'hab04: y = 16'hfe00;
			16'hab05: y = 16'hfe00;
			16'hab06: y = 16'hfe00;
			16'hab07: y = 16'hfe00;
			16'hab08: y = 16'hfe00;
			16'hab09: y = 16'hfe00;
			16'hab0a: y = 16'hfe00;
			16'hab0b: y = 16'hfe00;
			16'hab0c: y = 16'hfe00;
			16'hab0d: y = 16'hfe00;
			16'hab0e: y = 16'hfe00;
			16'hab0f: y = 16'hfe00;
			16'hab10: y = 16'hfe00;
			16'hab11: y = 16'hfe00;
			16'hab12: y = 16'hfe00;
			16'hab13: y = 16'hfe00;
			16'hab14: y = 16'hfe00;
			16'hab15: y = 16'hfe00;
			16'hab16: y = 16'hfe00;
			16'hab17: y = 16'hfe00;
			16'hab18: y = 16'hfe00;
			16'hab19: y = 16'hfe00;
			16'hab1a: y = 16'hfe00;
			16'hab1b: y = 16'hfe00;
			16'hab1c: y = 16'hfe00;
			16'hab1d: y = 16'hfe00;
			16'hab1e: y = 16'hfe00;
			16'hab1f: y = 16'hfe00;
			16'hab20: y = 16'hfe00;
			16'hab21: y = 16'hfe00;
			16'hab22: y = 16'hfe00;
			16'hab23: y = 16'hfe00;
			16'hab24: y = 16'hfe00;
			16'hab25: y = 16'hfe00;
			16'hab26: y = 16'hfe00;
			16'hab27: y = 16'hfe00;
			16'hab28: y = 16'hfe00;
			16'hab29: y = 16'hfe00;
			16'hab2a: y = 16'hfe00;
			16'hab2b: y = 16'hfe00;
			16'hab2c: y = 16'hfe00;
			16'hab2d: y = 16'hfe00;
			16'hab2e: y = 16'hfe00;
			16'hab2f: y = 16'hfe00;
			16'hab30: y = 16'hfe00;
			16'hab31: y = 16'hfe00;
			16'hab32: y = 16'hfe00;
			16'hab33: y = 16'hfe00;
			16'hab34: y = 16'hfe00;
			16'hab35: y = 16'hfe00;
			16'hab36: y = 16'hfe00;
			16'hab37: y = 16'hfe00;
			16'hab38: y = 16'hfe00;
			16'hab39: y = 16'hfe00;
			16'hab3a: y = 16'hfe00;
			16'hab3b: y = 16'hfe00;
			16'hab3c: y = 16'hfe00;
			16'hab3d: y = 16'hfe00;
			16'hab3e: y = 16'hfe00;
			16'hab3f: y = 16'hfe00;
			16'hab40: y = 16'hfe00;
			16'hab41: y = 16'hfe00;
			16'hab42: y = 16'hfe00;
			16'hab43: y = 16'hfe00;
			16'hab44: y = 16'hfe00;
			16'hab45: y = 16'hfe00;
			16'hab46: y = 16'hfe00;
			16'hab47: y = 16'hfe00;
			16'hab48: y = 16'hfe00;
			16'hab49: y = 16'hfe00;
			16'hab4a: y = 16'hfe00;
			16'hab4b: y = 16'hfe00;
			16'hab4c: y = 16'hfe00;
			16'hab4d: y = 16'hfe00;
			16'hab4e: y = 16'hfe00;
			16'hab4f: y = 16'hfe00;
			16'hab50: y = 16'hfe00;
			16'hab51: y = 16'hfe00;
			16'hab52: y = 16'hfe00;
			16'hab53: y = 16'hfe00;
			16'hab54: y = 16'hfe00;
			16'hab55: y = 16'hfe00;
			16'hab56: y = 16'hfe00;
			16'hab57: y = 16'hfe00;
			16'hab58: y = 16'hfe00;
			16'hab59: y = 16'hfe00;
			16'hab5a: y = 16'hfe00;
			16'hab5b: y = 16'hfe00;
			16'hab5c: y = 16'hfe00;
			16'hab5d: y = 16'hfe00;
			16'hab5e: y = 16'hfe00;
			16'hab5f: y = 16'hfe00;
			16'hab60: y = 16'hfe00;
			16'hab61: y = 16'hfe00;
			16'hab62: y = 16'hfe00;
			16'hab63: y = 16'hfe00;
			16'hab64: y = 16'hfe00;
			16'hab65: y = 16'hfe00;
			16'hab66: y = 16'hfe00;
			16'hab67: y = 16'hfe00;
			16'hab68: y = 16'hfe00;
			16'hab69: y = 16'hfe00;
			16'hab6a: y = 16'hfe00;
			16'hab6b: y = 16'hfe00;
			16'hab6c: y = 16'hfe00;
			16'hab6d: y = 16'hfe00;
			16'hab6e: y = 16'hfe00;
			16'hab6f: y = 16'hfe00;
			16'hab70: y = 16'hfe00;
			16'hab71: y = 16'hfe00;
			16'hab72: y = 16'hfe00;
			16'hab73: y = 16'hfe00;
			16'hab74: y = 16'hfe00;
			16'hab75: y = 16'hfe00;
			16'hab76: y = 16'hfe00;
			16'hab77: y = 16'hfe00;
			16'hab78: y = 16'hfe00;
			16'hab79: y = 16'hfe00;
			16'hab7a: y = 16'hfe00;
			16'hab7b: y = 16'hfe00;
			16'hab7c: y = 16'hfe00;
			16'hab7d: y = 16'hfe00;
			16'hab7e: y = 16'hfe00;
			16'hab7f: y = 16'hfe00;
			16'hab80: y = 16'hfe00;
			16'hab81: y = 16'hfe00;
			16'hab82: y = 16'hfe00;
			16'hab83: y = 16'hfe00;
			16'hab84: y = 16'hfe00;
			16'hab85: y = 16'hfe00;
			16'hab86: y = 16'hfe00;
			16'hab87: y = 16'hfe00;
			16'hab88: y = 16'hfe00;
			16'hab89: y = 16'hfe00;
			16'hab8a: y = 16'hfe00;
			16'hab8b: y = 16'hfe00;
			16'hab8c: y = 16'hfe00;
			16'hab8d: y = 16'hfe00;
			16'hab8e: y = 16'hfe00;
			16'hab8f: y = 16'hfe00;
			16'hab90: y = 16'hfe00;
			16'hab91: y = 16'hfe00;
			16'hab92: y = 16'hfe00;
			16'hab93: y = 16'hfe00;
			16'hab94: y = 16'hfe00;
			16'hab95: y = 16'hfe00;
			16'hab96: y = 16'hfe00;
			16'hab97: y = 16'hfe00;
			16'hab98: y = 16'hfe00;
			16'hab99: y = 16'hfe00;
			16'hab9a: y = 16'hfe00;
			16'hab9b: y = 16'hfe00;
			16'hab9c: y = 16'hfe00;
			16'hab9d: y = 16'hfe00;
			16'hab9e: y = 16'hfe00;
			16'hab9f: y = 16'hfe00;
			16'haba0: y = 16'hfe00;
			16'haba1: y = 16'hfe00;
			16'haba2: y = 16'hfe00;
			16'haba3: y = 16'hfe00;
			16'haba4: y = 16'hfe00;
			16'haba5: y = 16'hfe00;
			16'haba6: y = 16'hfe00;
			16'haba7: y = 16'hfe00;
			16'haba8: y = 16'hfe00;
			16'haba9: y = 16'hfe00;
			16'habaa: y = 16'hfe00;
			16'habab: y = 16'hfe00;
			16'habac: y = 16'hfe00;
			16'habad: y = 16'hfe00;
			16'habae: y = 16'hfe00;
			16'habaf: y = 16'hfe00;
			16'habb0: y = 16'hfe00;
			16'habb1: y = 16'hfe00;
			16'habb2: y = 16'hfe00;
			16'habb3: y = 16'hfe00;
			16'habb4: y = 16'hfe00;
			16'habb5: y = 16'hfe00;
			16'habb6: y = 16'hfe00;
			16'habb7: y = 16'hfe00;
			16'habb8: y = 16'hfe00;
			16'habb9: y = 16'hfe00;
			16'habba: y = 16'hfe00;
			16'habbb: y = 16'hfe00;
			16'habbc: y = 16'hfe00;
			16'habbd: y = 16'hfe00;
			16'habbe: y = 16'hfe00;
			16'habbf: y = 16'hfe00;
			16'habc0: y = 16'hfe00;
			16'habc1: y = 16'hfe00;
			16'habc2: y = 16'hfe00;
			16'habc3: y = 16'hfe00;
			16'habc4: y = 16'hfe00;
			16'habc5: y = 16'hfe00;
			16'habc6: y = 16'hfe00;
			16'habc7: y = 16'hfe00;
			16'habc8: y = 16'hfe00;
			16'habc9: y = 16'hfe00;
			16'habca: y = 16'hfe00;
			16'habcb: y = 16'hfe00;
			16'habcc: y = 16'hfe00;
			16'habcd: y = 16'hfe00;
			16'habce: y = 16'hfe00;
			16'habcf: y = 16'hfe00;
			16'habd0: y = 16'hfe00;
			16'habd1: y = 16'hfe00;
			16'habd2: y = 16'hfe00;
			16'habd3: y = 16'hfe00;
			16'habd4: y = 16'hfe00;
			16'habd5: y = 16'hfe00;
			16'habd6: y = 16'hfe00;
			16'habd7: y = 16'hfe00;
			16'habd8: y = 16'hfe00;
			16'habd9: y = 16'hfe00;
			16'habda: y = 16'hfe00;
			16'habdb: y = 16'hfe00;
			16'habdc: y = 16'hfe00;
			16'habdd: y = 16'hfe00;
			16'habde: y = 16'hfe00;
			16'habdf: y = 16'hfe00;
			16'habe0: y = 16'hfe00;
			16'habe1: y = 16'hfe00;
			16'habe2: y = 16'hfe00;
			16'habe3: y = 16'hfe00;
			16'habe4: y = 16'hfe00;
			16'habe5: y = 16'hfe00;
			16'habe6: y = 16'hfe00;
			16'habe7: y = 16'hfe00;
			16'habe8: y = 16'hfe00;
			16'habe9: y = 16'hfe00;
			16'habea: y = 16'hfe00;
			16'habeb: y = 16'hfe00;
			16'habec: y = 16'hfe00;
			16'habed: y = 16'hfe00;
			16'habee: y = 16'hfe00;
			16'habef: y = 16'hfe00;
			16'habf0: y = 16'hfe00;
			16'habf1: y = 16'hfe00;
			16'habf2: y = 16'hfe00;
			16'habf3: y = 16'hfe00;
			16'habf4: y = 16'hfe00;
			16'habf5: y = 16'hfe00;
			16'habf6: y = 16'hfe00;
			16'habf7: y = 16'hfe00;
			16'habf8: y = 16'hfe00;
			16'habf9: y = 16'hfe00;
			16'habfa: y = 16'hfe00;
			16'habfb: y = 16'hfe00;
			16'habfc: y = 16'hfe00;
			16'habfd: y = 16'hfe00;
			16'habfe: y = 16'hfe00;
			16'habff: y = 16'hfe00;
			16'hac00: y = 16'hfe00;
			16'hac01: y = 16'hfe00;
			16'hac02: y = 16'hfe00;
			16'hac03: y = 16'hfe00;
			16'hac04: y = 16'hfe00;
			16'hac05: y = 16'hfe00;
			16'hac06: y = 16'hfe00;
			16'hac07: y = 16'hfe00;
			16'hac08: y = 16'hfe00;
			16'hac09: y = 16'hfe00;
			16'hac0a: y = 16'hfe00;
			16'hac0b: y = 16'hfe00;
			16'hac0c: y = 16'hfe00;
			16'hac0d: y = 16'hfe00;
			16'hac0e: y = 16'hfe00;
			16'hac0f: y = 16'hfe00;
			16'hac10: y = 16'hfe00;
			16'hac11: y = 16'hfe00;
			16'hac12: y = 16'hfe00;
			16'hac13: y = 16'hfe00;
			16'hac14: y = 16'hfe00;
			16'hac15: y = 16'hfe00;
			16'hac16: y = 16'hfe00;
			16'hac17: y = 16'hfe00;
			16'hac18: y = 16'hfe00;
			16'hac19: y = 16'hfe00;
			16'hac1a: y = 16'hfe00;
			16'hac1b: y = 16'hfe00;
			16'hac1c: y = 16'hfe00;
			16'hac1d: y = 16'hfe00;
			16'hac1e: y = 16'hfe00;
			16'hac1f: y = 16'hfe00;
			16'hac20: y = 16'hfe00;
			16'hac21: y = 16'hfe00;
			16'hac22: y = 16'hfe00;
			16'hac23: y = 16'hfe00;
			16'hac24: y = 16'hfe00;
			16'hac25: y = 16'hfe00;
			16'hac26: y = 16'hfe00;
			16'hac27: y = 16'hfe00;
			16'hac28: y = 16'hfe00;
			16'hac29: y = 16'hfe00;
			16'hac2a: y = 16'hfe00;
			16'hac2b: y = 16'hfe00;
			16'hac2c: y = 16'hfe00;
			16'hac2d: y = 16'hfe00;
			16'hac2e: y = 16'hfe00;
			16'hac2f: y = 16'hfe00;
			16'hac30: y = 16'hfe00;
			16'hac31: y = 16'hfe00;
			16'hac32: y = 16'hfe00;
			16'hac33: y = 16'hfe00;
			16'hac34: y = 16'hfe00;
			16'hac35: y = 16'hfe00;
			16'hac36: y = 16'hfe00;
			16'hac37: y = 16'hfe00;
			16'hac38: y = 16'hfe00;
			16'hac39: y = 16'hfe00;
			16'hac3a: y = 16'hfe00;
			16'hac3b: y = 16'hfe00;
			16'hac3c: y = 16'hfe00;
			16'hac3d: y = 16'hfe00;
			16'hac3e: y = 16'hfe00;
			16'hac3f: y = 16'hfe00;
			16'hac40: y = 16'hfe00;
			16'hac41: y = 16'hfe00;
			16'hac42: y = 16'hfe00;
			16'hac43: y = 16'hfe00;
			16'hac44: y = 16'hfe00;
			16'hac45: y = 16'hfe00;
			16'hac46: y = 16'hfe00;
			16'hac47: y = 16'hfe00;
			16'hac48: y = 16'hfe00;
			16'hac49: y = 16'hfe00;
			16'hac4a: y = 16'hfe00;
			16'hac4b: y = 16'hfe00;
			16'hac4c: y = 16'hfe00;
			16'hac4d: y = 16'hfe00;
			16'hac4e: y = 16'hfe00;
			16'hac4f: y = 16'hfe00;
			16'hac50: y = 16'hfe00;
			16'hac51: y = 16'hfe00;
			16'hac52: y = 16'hfe00;
			16'hac53: y = 16'hfe00;
			16'hac54: y = 16'hfe00;
			16'hac55: y = 16'hfe00;
			16'hac56: y = 16'hfe00;
			16'hac57: y = 16'hfe00;
			16'hac58: y = 16'hfe00;
			16'hac59: y = 16'hfe00;
			16'hac5a: y = 16'hfe00;
			16'hac5b: y = 16'hfe00;
			16'hac5c: y = 16'hfe00;
			16'hac5d: y = 16'hfe00;
			16'hac5e: y = 16'hfe00;
			16'hac5f: y = 16'hfe00;
			16'hac60: y = 16'hfe00;
			16'hac61: y = 16'hfe00;
			16'hac62: y = 16'hfe00;
			16'hac63: y = 16'hfe00;
			16'hac64: y = 16'hfe00;
			16'hac65: y = 16'hfe00;
			16'hac66: y = 16'hfe00;
			16'hac67: y = 16'hfe00;
			16'hac68: y = 16'hfe00;
			16'hac69: y = 16'hfe00;
			16'hac6a: y = 16'hfe00;
			16'hac6b: y = 16'hfe00;
			16'hac6c: y = 16'hfe00;
			16'hac6d: y = 16'hfe00;
			16'hac6e: y = 16'hfe00;
			16'hac6f: y = 16'hfe00;
			16'hac70: y = 16'hfe00;
			16'hac71: y = 16'hfe00;
			16'hac72: y = 16'hfe00;
			16'hac73: y = 16'hfe00;
			16'hac74: y = 16'hfe00;
			16'hac75: y = 16'hfe00;
			16'hac76: y = 16'hfe00;
			16'hac77: y = 16'hfe00;
			16'hac78: y = 16'hfe00;
			16'hac79: y = 16'hfe00;
			16'hac7a: y = 16'hfe00;
			16'hac7b: y = 16'hfe00;
			16'hac7c: y = 16'hfe00;
			16'hac7d: y = 16'hfe00;
			16'hac7e: y = 16'hfe00;
			16'hac7f: y = 16'hfe00;
			16'hac80: y = 16'hfe00;
			16'hac81: y = 16'hfe00;
			16'hac82: y = 16'hfe00;
			16'hac83: y = 16'hfe00;
			16'hac84: y = 16'hfe00;
			16'hac85: y = 16'hfe00;
			16'hac86: y = 16'hfe00;
			16'hac87: y = 16'hfe00;
			16'hac88: y = 16'hfe00;
			16'hac89: y = 16'hfe00;
			16'hac8a: y = 16'hfe00;
			16'hac8b: y = 16'hfe00;
			16'hac8c: y = 16'hfe00;
			16'hac8d: y = 16'hfe00;
			16'hac8e: y = 16'hfe00;
			16'hac8f: y = 16'hfe00;
			16'hac90: y = 16'hfe00;
			16'hac91: y = 16'hfe00;
			16'hac92: y = 16'hfe00;
			16'hac93: y = 16'hfe00;
			16'hac94: y = 16'hfe00;
			16'hac95: y = 16'hfe00;
			16'hac96: y = 16'hfe00;
			16'hac97: y = 16'hfe00;
			16'hac98: y = 16'hfe00;
			16'hac99: y = 16'hfe00;
			16'hac9a: y = 16'hfe00;
			16'hac9b: y = 16'hfe00;
			16'hac9c: y = 16'hfe00;
			16'hac9d: y = 16'hfe00;
			16'hac9e: y = 16'hfe00;
			16'hac9f: y = 16'hfe00;
			16'haca0: y = 16'hfe00;
			16'haca1: y = 16'hfe00;
			16'haca2: y = 16'hfe00;
			16'haca3: y = 16'hfe00;
			16'haca4: y = 16'hfe00;
			16'haca5: y = 16'hfe00;
			16'haca6: y = 16'hfe00;
			16'haca7: y = 16'hfe00;
			16'haca8: y = 16'hfe00;
			16'haca9: y = 16'hfe00;
			16'hacaa: y = 16'hfe00;
			16'hacab: y = 16'hfe00;
			16'hacac: y = 16'hfe00;
			16'hacad: y = 16'hfe00;
			16'hacae: y = 16'hfe00;
			16'hacaf: y = 16'hfe00;
			16'hacb0: y = 16'hfe00;
			16'hacb1: y = 16'hfe00;
			16'hacb2: y = 16'hfe00;
			16'hacb3: y = 16'hfe00;
			16'hacb4: y = 16'hfe00;
			16'hacb5: y = 16'hfe00;
			16'hacb6: y = 16'hfe00;
			16'hacb7: y = 16'hfe00;
			16'hacb8: y = 16'hfe00;
			16'hacb9: y = 16'hfe00;
			16'hacba: y = 16'hfe00;
			16'hacbb: y = 16'hfe00;
			16'hacbc: y = 16'hfe00;
			16'hacbd: y = 16'hfe00;
			16'hacbe: y = 16'hfe00;
			16'hacbf: y = 16'hfe00;
			16'hacc0: y = 16'hfe00;
			16'hacc1: y = 16'hfe00;
			16'hacc2: y = 16'hfe00;
			16'hacc3: y = 16'hfe00;
			16'hacc4: y = 16'hfe00;
			16'hacc5: y = 16'hfe00;
			16'hacc6: y = 16'hfe00;
			16'hacc7: y = 16'hfe00;
			16'hacc8: y = 16'hfe00;
			16'hacc9: y = 16'hfe00;
			16'hacca: y = 16'hfe00;
			16'haccb: y = 16'hfe00;
			16'haccc: y = 16'hfe00;
			16'haccd: y = 16'hfe00;
			16'hacce: y = 16'hfe00;
			16'haccf: y = 16'hfe00;
			16'hacd0: y = 16'hfe00;
			16'hacd1: y = 16'hfe00;
			16'hacd2: y = 16'hfe00;
			16'hacd3: y = 16'hfe00;
			16'hacd4: y = 16'hfe00;
			16'hacd5: y = 16'hfe00;
			16'hacd6: y = 16'hfe00;
			16'hacd7: y = 16'hfe00;
			16'hacd8: y = 16'hfe00;
			16'hacd9: y = 16'hfe00;
			16'hacda: y = 16'hfe00;
			16'hacdb: y = 16'hfe00;
			16'hacdc: y = 16'hfe00;
			16'hacdd: y = 16'hfe00;
			16'hacde: y = 16'hfe00;
			16'hacdf: y = 16'hfe00;
			16'hace0: y = 16'hfe00;
			16'hace1: y = 16'hfe00;
			16'hace2: y = 16'hfe00;
			16'hace3: y = 16'hfe00;
			16'hace4: y = 16'hfe00;
			16'hace5: y = 16'hfe00;
			16'hace6: y = 16'hfe00;
			16'hace7: y = 16'hfe00;
			16'hace8: y = 16'hfe00;
			16'hace9: y = 16'hfe00;
			16'hacea: y = 16'hfe00;
			16'haceb: y = 16'hfe00;
			16'hacec: y = 16'hfe00;
			16'haced: y = 16'hfe00;
			16'hacee: y = 16'hfe00;
			16'hacef: y = 16'hfe00;
			16'hacf0: y = 16'hfe00;
			16'hacf1: y = 16'hfe00;
			16'hacf2: y = 16'hfe00;
			16'hacf3: y = 16'hfe00;
			16'hacf4: y = 16'hfe00;
			16'hacf5: y = 16'hfe00;
			16'hacf6: y = 16'hfe00;
			16'hacf7: y = 16'hfe00;
			16'hacf8: y = 16'hfe00;
			16'hacf9: y = 16'hfe00;
			16'hacfa: y = 16'hfe00;
			16'hacfb: y = 16'hfe00;
			16'hacfc: y = 16'hfe00;
			16'hacfd: y = 16'hfe00;
			16'hacfe: y = 16'hfe00;
			16'hacff: y = 16'hfe00;
			16'had00: y = 16'hfe00;
			16'had01: y = 16'hfe00;
			16'had02: y = 16'hfe00;
			16'had03: y = 16'hfe00;
			16'had04: y = 16'hfe00;
			16'had05: y = 16'hfe00;
			16'had06: y = 16'hfe00;
			16'had07: y = 16'hfe00;
			16'had08: y = 16'hfe00;
			16'had09: y = 16'hfe00;
			16'had0a: y = 16'hfe00;
			16'had0b: y = 16'hfe00;
			16'had0c: y = 16'hfe00;
			16'had0d: y = 16'hfe00;
			16'had0e: y = 16'hfe00;
			16'had0f: y = 16'hfe00;
			16'had10: y = 16'hfe00;
			16'had11: y = 16'hfe00;
			16'had12: y = 16'hfe00;
			16'had13: y = 16'hfe00;
			16'had14: y = 16'hfe00;
			16'had15: y = 16'hfe00;
			16'had16: y = 16'hfe00;
			16'had17: y = 16'hfe00;
			16'had18: y = 16'hfe00;
			16'had19: y = 16'hfe00;
			16'had1a: y = 16'hfe00;
			16'had1b: y = 16'hfe00;
			16'had1c: y = 16'hfe00;
			16'had1d: y = 16'hfe00;
			16'had1e: y = 16'hfe00;
			16'had1f: y = 16'hfe00;
			16'had20: y = 16'hfe00;
			16'had21: y = 16'hfe00;
			16'had22: y = 16'hfe00;
			16'had23: y = 16'hfe00;
			16'had24: y = 16'hfe00;
			16'had25: y = 16'hfe00;
			16'had26: y = 16'hfe00;
			16'had27: y = 16'hfe00;
			16'had28: y = 16'hfe00;
			16'had29: y = 16'hfe00;
			16'had2a: y = 16'hfe00;
			16'had2b: y = 16'hfe00;
			16'had2c: y = 16'hfe00;
			16'had2d: y = 16'hfe00;
			16'had2e: y = 16'hfe00;
			16'had2f: y = 16'hfe00;
			16'had30: y = 16'hfe00;
			16'had31: y = 16'hfe00;
			16'had32: y = 16'hfe00;
			16'had33: y = 16'hfe00;
			16'had34: y = 16'hfe00;
			16'had35: y = 16'hfe00;
			16'had36: y = 16'hfe00;
			16'had37: y = 16'hfe00;
			16'had38: y = 16'hfe00;
			16'had39: y = 16'hfe00;
			16'had3a: y = 16'hfe00;
			16'had3b: y = 16'hfe00;
			16'had3c: y = 16'hfe00;
			16'had3d: y = 16'hfe00;
			16'had3e: y = 16'hfe00;
			16'had3f: y = 16'hfe00;
			16'had40: y = 16'hfe00;
			16'had41: y = 16'hfe00;
			16'had42: y = 16'hfe00;
			16'had43: y = 16'hfe00;
			16'had44: y = 16'hfe00;
			16'had45: y = 16'hfe00;
			16'had46: y = 16'hfe00;
			16'had47: y = 16'hfe00;
			16'had48: y = 16'hfe00;
			16'had49: y = 16'hfe00;
			16'had4a: y = 16'hfe00;
			16'had4b: y = 16'hfe00;
			16'had4c: y = 16'hfe00;
			16'had4d: y = 16'hfe00;
			16'had4e: y = 16'hfe00;
			16'had4f: y = 16'hfe00;
			16'had50: y = 16'hfe00;
			16'had51: y = 16'hfe00;
			16'had52: y = 16'hfe00;
			16'had53: y = 16'hfe00;
			16'had54: y = 16'hfe00;
			16'had55: y = 16'hfe00;
			16'had56: y = 16'hfe00;
			16'had57: y = 16'hfe00;
			16'had58: y = 16'hfe00;
			16'had59: y = 16'hfe00;
			16'had5a: y = 16'hfe00;
			16'had5b: y = 16'hfe00;
			16'had5c: y = 16'hfe00;
			16'had5d: y = 16'hfe00;
			16'had5e: y = 16'hfe00;
			16'had5f: y = 16'hfe00;
			16'had60: y = 16'hfe00;
			16'had61: y = 16'hfe00;
			16'had62: y = 16'hfe00;
			16'had63: y = 16'hfe00;
			16'had64: y = 16'hfe00;
			16'had65: y = 16'hfe00;
			16'had66: y = 16'hfe00;
			16'had67: y = 16'hfe00;
			16'had68: y = 16'hfe00;
			16'had69: y = 16'hfe00;
			16'had6a: y = 16'hfe00;
			16'had6b: y = 16'hfe00;
			16'had6c: y = 16'hfe00;
			16'had6d: y = 16'hfe00;
			16'had6e: y = 16'hfe00;
			16'had6f: y = 16'hfe00;
			16'had70: y = 16'hfe00;
			16'had71: y = 16'hfe00;
			16'had72: y = 16'hfe00;
			16'had73: y = 16'hfe00;
			16'had74: y = 16'hfe00;
			16'had75: y = 16'hfe00;
			16'had76: y = 16'hfe00;
			16'had77: y = 16'hfe00;
			16'had78: y = 16'hfe00;
			16'had79: y = 16'hfe00;
			16'had7a: y = 16'hfe00;
			16'had7b: y = 16'hfe00;
			16'had7c: y = 16'hfe00;
			16'had7d: y = 16'hfe00;
			16'had7e: y = 16'hfe00;
			16'had7f: y = 16'hfe00;
			16'had80: y = 16'hfe00;
			16'had81: y = 16'hfe00;
			16'had82: y = 16'hfe00;
			16'had83: y = 16'hfe00;
			16'had84: y = 16'hfe00;
			16'had85: y = 16'hfe00;
			16'had86: y = 16'hfe00;
			16'had87: y = 16'hfe00;
			16'had88: y = 16'hfe00;
			16'had89: y = 16'hfe00;
			16'had8a: y = 16'hfe00;
			16'had8b: y = 16'hfe00;
			16'had8c: y = 16'hfe00;
			16'had8d: y = 16'hfe00;
			16'had8e: y = 16'hfe00;
			16'had8f: y = 16'hfe00;
			16'had90: y = 16'hfe00;
			16'had91: y = 16'hfe00;
			16'had92: y = 16'hfe00;
			16'had93: y = 16'hfe00;
			16'had94: y = 16'hfe00;
			16'had95: y = 16'hfe00;
			16'had96: y = 16'hfe00;
			16'had97: y = 16'hfe00;
			16'had98: y = 16'hfe00;
			16'had99: y = 16'hfe00;
			16'had9a: y = 16'hfe00;
			16'had9b: y = 16'hfe00;
			16'had9c: y = 16'hfe00;
			16'had9d: y = 16'hfe00;
			16'had9e: y = 16'hfe00;
			16'had9f: y = 16'hfe00;
			16'hada0: y = 16'hfe00;
			16'hada1: y = 16'hfe00;
			16'hada2: y = 16'hfe00;
			16'hada3: y = 16'hfe00;
			16'hada4: y = 16'hfe00;
			16'hada5: y = 16'hfe00;
			16'hada6: y = 16'hfe00;
			16'hada7: y = 16'hfe00;
			16'hada8: y = 16'hfe00;
			16'hada9: y = 16'hfe00;
			16'hadaa: y = 16'hfe00;
			16'hadab: y = 16'hfe00;
			16'hadac: y = 16'hfe00;
			16'hadad: y = 16'hfe00;
			16'hadae: y = 16'hfe00;
			16'hadaf: y = 16'hfe00;
			16'hadb0: y = 16'hfe00;
			16'hadb1: y = 16'hfe00;
			16'hadb2: y = 16'hfe00;
			16'hadb3: y = 16'hfe00;
			16'hadb4: y = 16'hfe00;
			16'hadb5: y = 16'hfe00;
			16'hadb6: y = 16'hfe00;
			16'hadb7: y = 16'hfe00;
			16'hadb8: y = 16'hfe00;
			16'hadb9: y = 16'hfe00;
			16'hadba: y = 16'hfe00;
			16'hadbb: y = 16'hfe00;
			16'hadbc: y = 16'hfe00;
			16'hadbd: y = 16'hfe00;
			16'hadbe: y = 16'hfe00;
			16'hadbf: y = 16'hfe00;
			16'hadc0: y = 16'hfe00;
			16'hadc1: y = 16'hfe00;
			16'hadc2: y = 16'hfe00;
			16'hadc3: y = 16'hfe00;
			16'hadc4: y = 16'hfe00;
			16'hadc5: y = 16'hfe00;
			16'hadc6: y = 16'hfe00;
			16'hadc7: y = 16'hfe00;
			16'hadc8: y = 16'hfe00;
			16'hadc9: y = 16'hfe00;
			16'hadca: y = 16'hfe00;
			16'hadcb: y = 16'hfe00;
			16'hadcc: y = 16'hfe00;
			16'hadcd: y = 16'hfe00;
			16'hadce: y = 16'hfe00;
			16'hadcf: y = 16'hfe00;
			16'hadd0: y = 16'hfe00;
			16'hadd1: y = 16'hfe00;
			16'hadd2: y = 16'hfe00;
			16'hadd3: y = 16'hfe00;
			16'hadd4: y = 16'hfe00;
			16'hadd5: y = 16'hfe00;
			16'hadd6: y = 16'hfe00;
			16'hadd7: y = 16'hfe00;
			16'hadd8: y = 16'hfe00;
			16'hadd9: y = 16'hfe00;
			16'hadda: y = 16'hfe00;
			16'haddb: y = 16'hfe00;
			16'haddc: y = 16'hfe00;
			16'haddd: y = 16'hfe00;
			16'hadde: y = 16'hfe00;
			16'haddf: y = 16'hfe00;
			16'hade0: y = 16'hfe00;
			16'hade1: y = 16'hfe00;
			16'hade2: y = 16'hfe00;
			16'hade3: y = 16'hfe00;
			16'hade4: y = 16'hfe00;
			16'hade5: y = 16'hfe00;
			16'hade6: y = 16'hfe00;
			16'hade7: y = 16'hfe00;
			16'hade8: y = 16'hfe00;
			16'hade9: y = 16'hfe00;
			16'hadea: y = 16'hfe00;
			16'hadeb: y = 16'hfe00;
			16'hadec: y = 16'hfe00;
			16'haded: y = 16'hfe00;
			16'hadee: y = 16'hfe00;
			16'hadef: y = 16'hfe00;
			16'hadf0: y = 16'hfe00;
			16'hadf1: y = 16'hfe00;
			16'hadf2: y = 16'hfe00;
			16'hadf3: y = 16'hfe00;
			16'hadf4: y = 16'hfe00;
			16'hadf5: y = 16'hfe00;
			16'hadf6: y = 16'hfe00;
			16'hadf7: y = 16'hfe00;
			16'hadf8: y = 16'hfe00;
			16'hadf9: y = 16'hfe00;
			16'hadfa: y = 16'hfe00;
			16'hadfb: y = 16'hfe00;
			16'hadfc: y = 16'hfe00;
			16'hadfd: y = 16'hfe00;
			16'hadfe: y = 16'hfe00;
			16'hadff: y = 16'hfe00;
			16'hae00: y = 16'hfe00;
			16'hae01: y = 16'hfe00;
			16'hae02: y = 16'hfe00;
			16'hae03: y = 16'hfe00;
			16'hae04: y = 16'hfe00;
			16'hae05: y = 16'hfe00;
			16'hae06: y = 16'hfe00;
			16'hae07: y = 16'hfe00;
			16'hae08: y = 16'hfe00;
			16'hae09: y = 16'hfe00;
			16'hae0a: y = 16'hfe00;
			16'hae0b: y = 16'hfe00;
			16'hae0c: y = 16'hfe00;
			16'hae0d: y = 16'hfe00;
			16'hae0e: y = 16'hfe00;
			16'hae0f: y = 16'hfe00;
			16'hae10: y = 16'hfe00;
			16'hae11: y = 16'hfe00;
			16'hae12: y = 16'hfe00;
			16'hae13: y = 16'hfe00;
			16'hae14: y = 16'hfe00;
			16'hae15: y = 16'hfe00;
			16'hae16: y = 16'hfe00;
			16'hae17: y = 16'hfe00;
			16'hae18: y = 16'hfe00;
			16'hae19: y = 16'hfe00;
			16'hae1a: y = 16'hfe00;
			16'hae1b: y = 16'hfe00;
			16'hae1c: y = 16'hfe00;
			16'hae1d: y = 16'hfe00;
			16'hae1e: y = 16'hfe00;
			16'hae1f: y = 16'hfe00;
			16'hae20: y = 16'hfe00;
			16'hae21: y = 16'hfe00;
			16'hae22: y = 16'hfe00;
			16'hae23: y = 16'hfe00;
			16'hae24: y = 16'hfe00;
			16'hae25: y = 16'hfe00;
			16'hae26: y = 16'hfe00;
			16'hae27: y = 16'hfe00;
			16'hae28: y = 16'hfe00;
			16'hae29: y = 16'hfe00;
			16'hae2a: y = 16'hfe00;
			16'hae2b: y = 16'hfe00;
			16'hae2c: y = 16'hfe00;
			16'hae2d: y = 16'hfe00;
			16'hae2e: y = 16'hfe00;
			16'hae2f: y = 16'hfe00;
			16'hae30: y = 16'hfe00;
			16'hae31: y = 16'hfe00;
			16'hae32: y = 16'hfe00;
			16'hae33: y = 16'hfe00;
			16'hae34: y = 16'hfe00;
			16'hae35: y = 16'hfe00;
			16'hae36: y = 16'hfe00;
			16'hae37: y = 16'hfe00;
			16'hae38: y = 16'hfe00;
			16'hae39: y = 16'hfe00;
			16'hae3a: y = 16'hfe00;
			16'hae3b: y = 16'hfe00;
			16'hae3c: y = 16'hfe00;
			16'hae3d: y = 16'hfe00;
			16'hae3e: y = 16'hfe00;
			16'hae3f: y = 16'hfe00;
			16'hae40: y = 16'hfe00;
			16'hae41: y = 16'hfe00;
			16'hae42: y = 16'hfe00;
			16'hae43: y = 16'hfe00;
			16'hae44: y = 16'hfe00;
			16'hae45: y = 16'hfe00;
			16'hae46: y = 16'hfe00;
			16'hae47: y = 16'hfe00;
			16'hae48: y = 16'hfe00;
			16'hae49: y = 16'hfe00;
			16'hae4a: y = 16'hfe00;
			16'hae4b: y = 16'hfe00;
			16'hae4c: y = 16'hfe00;
			16'hae4d: y = 16'hfe00;
			16'hae4e: y = 16'hfe00;
			16'hae4f: y = 16'hfe00;
			16'hae50: y = 16'hfe00;
			16'hae51: y = 16'hfe00;
			16'hae52: y = 16'hfe00;
			16'hae53: y = 16'hfe00;
			16'hae54: y = 16'hfe00;
			16'hae55: y = 16'hfe00;
			16'hae56: y = 16'hfe00;
			16'hae57: y = 16'hfe00;
			16'hae58: y = 16'hfe00;
			16'hae59: y = 16'hfe00;
			16'hae5a: y = 16'hfe00;
			16'hae5b: y = 16'hfe00;
			16'hae5c: y = 16'hfe00;
			16'hae5d: y = 16'hfe00;
			16'hae5e: y = 16'hfe00;
			16'hae5f: y = 16'hfe00;
			16'hae60: y = 16'hfe00;
			16'hae61: y = 16'hfe00;
			16'hae62: y = 16'hfe00;
			16'hae63: y = 16'hfe00;
			16'hae64: y = 16'hfe00;
			16'hae65: y = 16'hfe00;
			16'hae66: y = 16'hfe00;
			16'hae67: y = 16'hfe00;
			16'hae68: y = 16'hfe00;
			16'hae69: y = 16'hfe00;
			16'hae6a: y = 16'hfe00;
			16'hae6b: y = 16'hfe00;
			16'hae6c: y = 16'hfe00;
			16'hae6d: y = 16'hfe00;
			16'hae6e: y = 16'hfe00;
			16'hae6f: y = 16'hfe00;
			16'hae70: y = 16'hfe00;
			16'hae71: y = 16'hfe00;
			16'hae72: y = 16'hfe00;
			16'hae73: y = 16'hfe00;
			16'hae74: y = 16'hfe00;
			16'hae75: y = 16'hfe00;
			16'hae76: y = 16'hfe00;
			16'hae77: y = 16'hfe00;
			16'hae78: y = 16'hfe00;
			16'hae79: y = 16'hfe00;
			16'hae7a: y = 16'hfe00;
			16'hae7b: y = 16'hfe00;
			16'hae7c: y = 16'hfe00;
			16'hae7d: y = 16'hfe00;
			16'hae7e: y = 16'hfe00;
			16'hae7f: y = 16'hfe00;
			16'hae80: y = 16'hfe00;
			16'hae81: y = 16'hfe00;
			16'hae82: y = 16'hfe00;
			16'hae83: y = 16'hfe00;
			16'hae84: y = 16'hfe00;
			16'hae85: y = 16'hfe00;
			16'hae86: y = 16'hfe00;
			16'hae87: y = 16'hfe00;
			16'hae88: y = 16'hfe00;
			16'hae89: y = 16'hfe00;
			16'hae8a: y = 16'hfe00;
			16'hae8b: y = 16'hfe00;
			16'hae8c: y = 16'hfe00;
			16'hae8d: y = 16'hfe00;
			16'hae8e: y = 16'hfe00;
			16'hae8f: y = 16'hfe00;
			16'hae90: y = 16'hfe00;
			16'hae91: y = 16'hfe00;
			16'hae92: y = 16'hfe00;
			16'hae93: y = 16'hfe00;
			16'hae94: y = 16'hfe00;
			16'hae95: y = 16'hfe00;
			16'hae96: y = 16'hfe00;
			16'hae97: y = 16'hfe00;
			16'hae98: y = 16'hfe00;
			16'hae99: y = 16'hfe00;
			16'hae9a: y = 16'hfe00;
			16'hae9b: y = 16'hfe00;
			16'hae9c: y = 16'hfe00;
			16'hae9d: y = 16'hfe00;
			16'hae9e: y = 16'hfe00;
			16'hae9f: y = 16'hfe00;
			16'haea0: y = 16'hfe00;
			16'haea1: y = 16'hfe00;
			16'haea2: y = 16'hfe00;
			16'haea3: y = 16'hfe00;
			16'haea4: y = 16'hfe00;
			16'haea5: y = 16'hfe00;
			16'haea6: y = 16'hfe00;
			16'haea7: y = 16'hfe00;
			16'haea8: y = 16'hfe00;
			16'haea9: y = 16'hfe00;
			16'haeaa: y = 16'hfe00;
			16'haeab: y = 16'hfe00;
			16'haeac: y = 16'hfe00;
			16'haead: y = 16'hfe00;
			16'haeae: y = 16'hfe00;
			16'haeaf: y = 16'hfe00;
			16'haeb0: y = 16'hfe00;
			16'haeb1: y = 16'hfe00;
			16'haeb2: y = 16'hfe00;
			16'haeb3: y = 16'hfe00;
			16'haeb4: y = 16'hfe00;
			16'haeb5: y = 16'hfe00;
			16'haeb6: y = 16'hfe00;
			16'haeb7: y = 16'hfe00;
			16'haeb8: y = 16'hfe00;
			16'haeb9: y = 16'hfe00;
			16'haeba: y = 16'hfe00;
			16'haebb: y = 16'hfe00;
			16'haebc: y = 16'hfe00;
			16'haebd: y = 16'hfe00;
			16'haebe: y = 16'hfe00;
			16'haebf: y = 16'hfe00;
			16'haec0: y = 16'hfe00;
			16'haec1: y = 16'hfe00;
			16'haec2: y = 16'hfe00;
			16'haec3: y = 16'hfe00;
			16'haec4: y = 16'hfe00;
			16'haec5: y = 16'hfe00;
			16'haec6: y = 16'hfe00;
			16'haec7: y = 16'hfe00;
			16'haec8: y = 16'hfe00;
			16'haec9: y = 16'hfe00;
			16'haeca: y = 16'hfe00;
			16'haecb: y = 16'hfe00;
			16'haecc: y = 16'hfe00;
			16'haecd: y = 16'hfe00;
			16'haece: y = 16'hfe00;
			16'haecf: y = 16'hfe00;
			16'haed0: y = 16'hfe00;
			16'haed1: y = 16'hfe00;
			16'haed2: y = 16'hfe00;
			16'haed3: y = 16'hfe00;
			16'haed4: y = 16'hfe00;
			16'haed5: y = 16'hfe00;
			16'haed6: y = 16'hfe00;
			16'haed7: y = 16'hfe00;
			16'haed8: y = 16'hfe00;
			16'haed9: y = 16'hfe00;
			16'haeda: y = 16'hfe00;
			16'haedb: y = 16'hfe00;
			16'haedc: y = 16'hfe00;
			16'haedd: y = 16'hfe00;
			16'haede: y = 16'hfe00;
			16'haedf: y = 16'hfe00;
			16'haee0: y = 16'hfe00;
			16'haee1: y = 16'hfe00;
			16'haee2: y = 16'hfe00;
			16'haee3: y = 16'hfe00;
			16'haee4: y = 16'hfe00;
			16'haee5: y = 16'hfe00;
			16'haee6: y = 16'hfe00;
			16'haee7: y = 16'hfe00;
			16'haee8: y = 16'hfe00;
			16'haee9: y = 16'hfe00;
			16'haeea: y = 16'hfe00;
			16'haeeb: y = 16'hfe00;
			16'haeec: y = 16'hfe00;
			16'haeed: y = 16'hfe00;
			16'haeee: y = 16'hfe00;
			16'haeef: y = 16'hfe00;
			16'haef0: y = 16'hfe00;
			16'haef1: y = 16'hfe00;
			16'haef2: y = 16'hfe00;
			16'haef3: y = 16'hfe00;
			16'haef4: y = 16'hfe00;
			16'haef5: y = 16'hfe00;
			16'haef6: y = 16'hfe00;
			16'haef7: y = 16'hfe00;
			16'haef8: y = 16'hfe00;
			16'haef9: y = 16'hfe00;
			16'haefa: y = 16'hfe00;
			16'haefb: y = 16'hfe00;
			16'haefc: y = 16'hfe00;
			16'haefd: y = 16'hfe00;
			16'haefe: y = 16'hfe00;
			16'haeff: y = 16'hfe00;
			16'haf00: y = 16'hfe00;
			16'haf01: y = 16'hfe00;
			16'haf02: y = 16'hfe00;
			16'haf03: y = 16'hfe00;
			16'haf04: y = 16'hfe00;
			16'haf05: y = 16'hfe00;
			16'haf06: y = 16'hfe00;
			16'haf07: y = 16'hfe00;
			16'haf08: y = 16'hfe00;
			16'haf09: y = 16'hfe00;
			16'haf0a: y = 16'hfe00;
			16'haf0b: y = 16'hfe00;
			16'haf0c: y = 16'hfe00;
			16'haf0d: y = 16'hfe00;
			16'haf0e: y = 16'hfe00;
			16'haf0f: y = 16'hfe00;
			16'haf10: y = 16'hfe00;
			16'haf11: y = 16'hfe00;
			16'haf12: y = 16'hfe00;
			16'haf13: y = 16'hfe00;
			16'haf14: y = 16'hfe00;
			16'haf15: y = 16'hfe00;
			16'haf16: y = 16'hfe00;
			16'haf17: y = 16'hfe00;
			16'haf18: y = 16'hfe00;
			16'haf19: y = 16'hfe00;
			16'haf1a: y = 16'hfe00;
			16'haf1b: y = 16'hfe00;
			16'haf1c: y = 16'hfe00;
			16'haf1d: y = 16'hfe00;
			16'haf1e: y = 16'hfe00;
			16'haf1f: y = 16'hfe00;
			16'haf20: y = 16'hfe00;
			16'haf21: y = 16'hfe00;
			16'haf22: y = 16'hfe00;
			16'haf23: y = 16'hfe00;
			16'haf24: y = 16'hfe00;
			16'haf25: y = 16'hfe00;
			16'haf26: y = 16'hfe00;
			16'haf27: y = 16'hfe00;
			16'haf28: y = 16'hfe00;
			16'haf29: y = 16'hfe00;
			16'haf2a: y = 16'hfe00;
			16'haf2b: y = 16'hfe00;
			16'haf2c: y = 16'hfe00;
			16'haf2d: y = 16'hfe00;
			16'haf2e: y = 16'hfe00;
			16'haf2f: y = 16'hfe00;
			16'haf30: y = 16'hfe00;
			16'haf31: y = 16'hfe00;
			16'haf32: y = 16'hfe00;
			16'haf33: y = 16'hfe00;
			16'haf34: y = 16'hfe00;
			16'haf35: y = 16'hfe00;
			16'haf36: y = 16'hfe00;
			16'haf37: y = 16'hfe00;
			16'haf38: y = 16'hfe00;
			16'haf39: y = 16'hfe00;
			16'haf3a: y = 16'hfe00;
			16'haf3b: y = 16'hfe00;
			16'haf3c: y = 16'hfe00;
			16'haf3d: y = 16'hfe00;
			16'haf3e: y = 16'hfe00;
			16'haf3f: y = 16'hfe00;
			16'haf40: y = 16'hfe00;
			16'haf41: y = 16'hfe00;
			16'haf42: y = 16'hfe00;
			16'haf43: y = 16'hfe00;
			16'haf44: y = 16'hfe00;
			16'haf45: y = 16'hfe00;
			16'haf46: y = 16'hfe00;
			16'haf47: y = 16'hfe00;
			16'haf48: y = 16'hfe00;
			16'haf49: y = 16'hfe00;
			16'haf4a: y = 16'hfe00;
			16'haf4b: y = 16'hfe00;
			16'haf4c: y = 16'hfe00;
			16'haf4d: y = 16'hfe00;
			16'haf4e: y = 16'hfe00;
			16'haf4f: y = 16'hfe00;
			16'haf50: y = 16'hfe00;
			16'haf51: y = 16'hfe00;
			16'haf52: y = 16'hfe00;
			16'haf53: y = 16'hfe00;
			16'haf54: y = 16'hfe00;
			16'haf55: y = 16'hfe00;
			16'haf56: y = 16'hfe00;
			16'haf57: y = 16'hfe00;
			16'haf58: y = 16'hfe00;
			16'haf59: y = 16'hfe00;
			16'haf5a: y = 16'hfe00;
			16'haf5b: y = 16'hfe00;
			16'haf5c: y = 16'hfe00;
			16'haf5d: y = 16'hfe00;
			16'haf5e: y = 16'hfe00;
			16'haf5f: y = 16'hfe00;
			16'haf60: y = 16'hfe00;
			16'haf61: y = 16'hfe00;
			16'haf62: y = 16'hfe00;
			16'haf63: y = 16'hfe00;
			16'haf64: y = 16'hfe00;
			16'haf65: y = 16'hfe00;
			16'haf66: y = 16'hfe00;
			16'haf67: y = 16'hfe00;
			16'haf68: y = 16'hfe00;
			16'haf69: y = 16'hfe00;
			16'haf6a: y = 16'hfe00;
			16'haf6b: y = 16'hfe00;
			16'haf6c: y = 16'hfe00;
			16'haf6d: y = 16'hfe00;
			16'haf6e: y = 16'hfe00;
			16'haf6f: y = 16'hfe00;
			16'haf70: y = 16'hfe00;
			16'haf71: y = 16'hfe00;
			16'haf72: y = 16'hfe00;
			16'haf73: y = 16'hfe00;
			16'haf74: y = 16'hfe00;
			16'haf75: y = 16'hfe00;
			16'haf76: y = 16'hfe00;
			16'haf77: y = 16'hfe00;
			16'haf78: y = 16'hfe00;
			16'haf79: y = 16'hfe00;
			16'haf7a: y = 16'hfe00;
			16'haf7b: y = 16'hfe00;
			16'haf7c: y = 16'hfe00;
			16'haf7d: y = 16'hfe00;
			16'haf7e: y = 16'hfe00;
			16'haf7f: y = 16'hfe00;
			16'haf80: y = 16'hfe00;
			16'haf81: y = 16'hfe00;
			16'haf82: y = 16'hfe00;
			16'haf83: y = 16'hfe00;
			16'haf84: y = 16'hfe00;
			16'haf85: y = 16'hfe00;
			16'haf86: y = 16'hfe00;
			16'haf87: y = 16'hfe00;
			16'haf88: y = 16'hfe00;
			16'haf89: y = 16'hfe00;
			16'haf8a: y = 16'hfe00;
			16'haf8b: y = 16'hfe00;
			16'haf8c: y = 16'hfe00;
			16'haf8d: y = 16'hfe00;
			16'haf8e: y = 16'hfe00;
			16'haf8f: y = 16'hfe00;
			16'haf90: y = 16'hfe00;
			16'haf91: y = 16'hfe00;
			16'haf92: y = 16'hfe00;
			16'haf93: y = 16'hfe00;
			16'haf94: y = 16'hfe00;
			16'haf95: y = 16'hfe00;
			16'haf96: y = 16'hfe00;
			16'haf97: y = 16'hfe00;
			16'haf98: y = 16'hfe00;
			16'haf99: y = 16'hfe00;
			16'haf9a: y = 16'hfe00;
			16'haf9b: y = 16'hfe00;
			16'haf9c: y = 16'hfe00;
			16'haf9d: y = 16'hfe00;
			16'haf9e: y = 16'hfe00;
			16'haf9f: y = 16'hfe00;
			16'hafa0: y = 16'hfe00;
			16'hafa1: y = 16'hfe00;
			16'hafa2: y = 16'hfe00;
			16'hafa3: y = 16'hfe00;
			16'hafa4: y = 16'hfe00;
			16'hafa5: y = 16'hfe00;
			16'hafa6: y = 16'hfe00;
			16'hafa7: y = 16'hfe00;
			16'hafa8: y = 16'hfe00;
			16'hafa9: y = 16'hfe00;
			16'hafaa: y = 16'hfe00;
			16'hafab: y = 16'hfe00;
			16'hafac: y = 16'hfe00;
			16'hafad: y = 16'hfe00;
			16'hafae: y = 16'hfe00;
			16'hafaf: y = 16'hfe00;
			16'hafb0: y = 16'hfe00;
			16'hafb1: y = 16'hfe00;
			16'hafb2: y = 16'hfe00;
			16'hafb3: y = 16'hfe00;
			16'hafb4: y = 16'hfe00;
			16'hafb5: y = 16'hfe00;
			16'hafb6: y = 16'hfe00;
			16'hafb7: y = 16'hfe00;
			16'hafb8: y = 16'hfe00;
			16'hafb9: y = 16'hfe00;
			16'hafba: y = 16'hfe00;
			16'hafbb: y = 16'hfe00;
			16'hafbc: y = 16'hfe00;
			16'hafbd: y = 16'hfe00;
			16'hafbe: y = 16'hfe00;
			16'hafbf: y = 16'hfe00;
			16'hafc0: y = 16'hfe00;
			16'hafc1: y = 16'hfe00;
			16'hafc2: y = 16'hfe00;
			16'hafc3: y = 16'hfe00;
			16'hafc4: y = 16'hfe00;
			16'hafc5: y = 16'hfe00;
			16'hafc6: y = 16'hfe00;
			16'hafc7: y = 16'hfe00;
			16'hafc8: y = 16'hfe00;
			16'hafc9: y = 16'hfe00;
			16'hafca: y = 16'hfe00;
			16'hafcb: y = 16'hfe00;
			16'hafcc: y = 16'hfe00;
			16'hafcd: y = 16'hfe00;
			16'hafce: y = 16'hfe00;
			16'hafcf: y = 16'hfe00;
			16'hafd0: y = 16'hfe00;
			16'hafd1: y = 16'hfe00;
			16'hafd2: y = 16'hfe00;
			16'hafd3: y = 16'hfe00;
			16'hafd4: y = 16'hfe00;
			16'hafd5: y = 16'hfe00;
			16'hafd6: y = 16'hfe00;
			16'hafd7: y = 16'hfe00;
			16'hafd8: y = 16'hfe00;
			16'hafd9: y = 16'hfe00;
			16'hafda: y = 16'hfe00;
			16'hafdb: y = 16'hfe00;
			16'hafdc: y = 16'hfe00;
			16'hafdd: y = 16'hfe00;
			16'hafde: y = 16'hfe00;
			16'hafdf: y = 16'hfe00;
			16'hafe0: y = 16'hfe00;
			16'hafe1: y = 16'hfe00;
			16'hafe2: y = 16'hfe00;
			16'hafe3: y = 16'hfe00;
			16'hafe4: y = 16'hfe00;
			16'hafe5: y = 16'hfe00;
			16'hafe6: y = 16'hfe00;
			16'hafe7: y = 16'hfe00;
			16'hafe8: y = 16'hfe00;
			16'hafe9: y = 16'hfe00;
			16'hafea: y = 16'hfe00;
			16'hafeb: y = 16'hfe00;
			16'hafec: y = 16'hfe00;
			16'hafed: y = 16'hfe00;
			16'hafee: y = 16'hfe00;
			16'hafef: y = 16'hfe00;
			16'haff0: y = 16'hfe00;
			16'haff1: y = 16'hfe00;
			16'haff2: y = 16'hfe00;
			16'haff3: y = 16'hfe00;
			16'haff4: y = 16'hfe00;
			16'haff5: y = 16'hfe00;
			16'haff6: y = 16'hfe00;
			16'haff7: y = 16'hfe00;
			16'haff8: y = 16'hfe00;
			16'haff9: y = 16'hfe00;
			16'haffa: y = 16'hfe00;
			16'haffb: y = 16'hfe00;
			16'haffc: y = 16'hfe00;
			16'haffd: y = 16'hfe00;
			16'haffe: y = 16'hfe00;
			16'hafff: y = 16'hfe00;
			16'hb000: y = 16'hfe00;
			16'hb001: y = 16'hfe00;
			16'hb002: y = 16'hfe00;
			16'hb003: y = 16'hfe00;
			16'hb004: y = 16'hfe00;
			16'hb005: y = 16'hfe00;
			16'hb006: y = 16'hfe00;
			16'hb007: y = 16'hfe00;
			16'hb008: y = 16'hfe00;
			16'hb009: y = 16'hfe00;
			16'hb00a: y = 16'hfe00;
			16'hb00b: y = 16'hfe00;
			16'hb00c: y = 16'hfe00;
			16'hb00d: y = 16'hfe00;
			16'hb00e: y = 16'hfe00;
			16'hb00f: y = 16'hfe00;
			16'hb010: y = 16'hfe00;
			16'hb011: y = 16'hfe00;
			16'hb012: y = 16'hfe00;
			16'hb013: y = 16'hfe00;
			16'hb014: y = 16'hfe00;
			16'hb015: y = 16'hfe00;
			16'hb016: y = 16'hfe00;
			16'hb017: y = 16'hfe00;
			16'hb018: y = 16'hfe00;
			16'hb019: y = 16'hfe00;
			16'hb01a: y = 16'hfe00;
			16'hb01b: y = 16'hfe00;
			16'hb01c: y = 16'hfe00;
			16'hb01d: y = 16'hfe00;
			16'hb01e: y = 16'hfe00;
			16'hb01f: y = 16'hfe00;
			16'hb020: y = 16'hfe00;
			16'hb021: y = 16'hfe00;
			16'hb022: y = 16'hfe00;
			16'hb023: y = 16'hfe00;
			16'hb024: y = 16'hfe00;
			16'hb025: y = 16'hfe00;
			16'hb026: y = 16'hfe00;
			16'hb027: y = 16'hfe00;
			16'hb028: y = 16'hfe00;
			16'hb029: y = 16'hfe00;
			16'hb02a: y = 16'hfe00;
			16'hb02b: y = 16'hfe00;
			16'hb02c: y = 16'hfe00;
			16'hb02d: y = 16'hfe00;
			16'hb02e: y = 16'hfe00;
			16'hb02f: y = 16'hfe00;
			16'hb030: y = 16'hfe00;
			16'hb031: y = 16'hfe00;
			16'hb032: y = 16'hfe00;
			16'hb033: y = 16'hfe00;
			16'hb034: y = 16'hfe00;
			16'hb035: y = 16'hfe00;
			16'hb036: y = 16'hfe00;
			16'hb037: y = 16'hfe00;
			16'hb038: y = 16'hfe00;
			16'hb039: y = 16'hfe00;
			16'hb03a: y = 16'hfe00;
			16'hb03b: y = 16'hfe00;
			16'hb03c: y = 16'hfe00;
			16'hb03d: y = 16'hfe00;
			16'hb03e: y = 16'hfe00;
			16'hb03f: y = 16'hfe00;
			16'hb040: y = 16'hfe00;
			16'hb041: y = 16'hfe00;
			16'hb042: y = 16'hfe00;
			16'hb043: y = 16'hfe00;
			16'hb044: y = 16'hfe00;
			16'hb045: y = 16'hfe00;
			16'hb046: y = 16'hfe00;
			16'hb047: y = 16'hfe00;
			16'hb048: y = 16'hfe00;
			16'hb049: y = 16'hfe00;
			16'hb04a: y = 16'hfe00;
			16'hb04b: y = 16'hfe00;
			16'hb04c: y = 16'hfe00;
			16'hb04d: y = 16'hfe00;
			16'hb04e: y = 16'hfe00;
			16'hb04f: y = 16'hfe00;
			16'hb050: y = 16'hfe00;
			16'hb051: y = 16'hfe00;
			16'hb052: y = 16'hfe00;
			16'hb053: y = 16'hfe00;
			16'hb054: y = 16'hfe00;
			16'hb055: y = 16'hfe00;
			16'hb056: y = 16'hfe00;
			16'hb057: y = 16'hfe00;
			16'hb058: y = 16'hfe00;
			16'hb059: y = 16'hfe00;
			16'hb05a: y = 16'hfe00;
			16'hb05b: y = 16'hfe00;
			16'hb05c: y = 16'hfe00;
			16'hb05d: y = 16'hfe00;
			16'hb05e: y = 16'hfe00;
			16'hb05f: y = 16'hfe00;
			16'hb060: y = 16'hfe00;
			16'hb061: y = 16'hfe00;
			16'hb062: y = 16'hfe00;
			16'hb063: y = 16'hfe00;
			16'hb064: y = 16'hfe00;
			16'hb065: y = 16'hfe00;
			16'hb066: y = 16'hfe00;
			16'hb067: y = 16'hfe00;
			16'hb068: y = 16'hfe00;
			16'hb069: y = 16'hfe00;
			16'hb06a: y = 16'hfe00;
			16'hb06b: y = 16'hfe00;
			16'hb06c: y = 16'hfe00;
			16'hb06d: y = 16'hfe00;
			16'hb06e: y = 16'hfe00;
			16'hb06f: y = 16'hfe00;
			16'hb070: y = 16'hfe00;
			16'hb071: y = 16'hfe00;
			16'hb072: y = 16'hfe00;
			16'hb073: y = 16'hfe00;
			16'hb074: y = 16'hfe00;
			16'hb075: y = 16'hfe00;
			16'hb076: y = 16'hfe00;
			16'hb077: y = 16'hfe00;
			16'hb078: y = 16'hfe00;
			16'hb079: y = 16'hfe00;
			16'hb07a: y = 16'hfe00;
			16'hb07b: y = 16'hfe00;
			16'hb07c: y = 16'hfe00;
			16'hb07d: y = 16'hfe00;
			16'hb07e: y = 16'hfe00;
			16'hb07f: y = 16'hfe00;
			16'hb080: y = 16'hfe00;
			16'hb081: y = 16'hfe00;
			16'hb082: y = 16'hfe00;
			16'hb083: y = 16'hfe00;
			16'hb084: y = 16'hfe00;
			16'hb085: y = 16'hfe00;
			16'hb086: y = 16'hfe00;
			16'hb087: y = 16'hfe00;
			16'hb088: y = 16'hfe00;
			16'hb089: y = 16'hfe00;
			16'hb08a: y = 16'hfe00;
			16'hb08b: y = 16'hfe00;
			16'hb08c: y = 16'hfe00;
			16'hb08d: y = 16'hfe00;
			16'hb08e: y = 16'hfe00;
			16'hb08f: y = 16'hfe00;
			16'hb090: y = 16'hfe00;
			16'hb091: y = 16'hfe00;
			16'hb092: y = 16'hfe00;
			16'hb093: y = 16'hfe00;
			16'hb094: y = 16'hfe00;
			16'hb095: y = 16'hfe00;
			16'hb096: y = 16'hfe00;
			16'hb097: y = 16'hfe00;
			16'hb098: y = 16'hfe00;
			16'hb099: y = 16'hfe00;
			16'hb09a: y = 16'hfe00;
			16'hb09b: y = 16'hfe00;
			16'hb09c: y = 16'hfe00;
			16'hb09d: y = 16'hfe00;
			16'hb09e: y = 16'hfe00;
			16'hb09f: y = 16'hfe00;
			16'hb0a0: y = 16'hfe00;
			16'hb0a1: y = 16'hfe00;
			16'hb0a2: y = 16'hfe00;
			16'hb0a3: y = 16'hfe00;
			16'hb0a4: y = 16'hfe00;
			16'hb0a5: y = 16'hfe00;
			16'hb0a6: y = 16'hfe00;
			16'hb0a7: y = 16'hfe00;
			16'hb0a8: y = 16'hfe00;
			16'hb0a9: y = 16'hfe00;
			16'hb0aa: y = 16'hfe00;
			16'hb0ab: y = 16'hfe00;
			16'hb0ac: y = 16'hfe00;
			16'hb0ad: y = 16'hfe00;
			16'hb0ae: y = 16'hfe00;
			16'hb0af: y = 16'hfe00;
			16'hb0b0: y = 16'hfe00;
			16'hb0b1: y = 16'hfe00;
			16'hb0b2: y = 16'hfe00;
			16'hb0b3: y = 16'hfe00;
			16'hb0b4: y = 16'hfe00;
			16'hb0b5: y = 16'hfe00;
			16'hb0b6: y = 16'hfe00;
			16'hb0b7: y = 16'hfe00;
			16'hb0b8: y = 16'hfe00;
			16'hb0b9: y = 16'hfe00;
			16'hb0ba: y = 16'hfe00;
			16'hb0bb: y = 16'hfe00;
			16'hb0bc: y = 16'hfe00;
			16'hb0bd: y = 16'hfe00;
			16'hb0be: y = 16'hfe00;
			16'hb0bf: y = 16'hfe00;
			16'hb0c0: y = 16'hfe00;
			16'hb0c1: y = 16'hfe00;
			16'hb0c2: y = 16'hfe00;
			16'hb0c3: y = 16'hfe00;
			16'hb0c4: y = 16'hfe00;
			16'hb0c5: y = 16'hfe00;
			16'hb0c6: y = 16'hfe00;
			16'hb0c7: y = 16'hfe00;
			16'hb0c8: y = 16'hfe00;
			16'hb0c9: y = 16'hfe00;
			16'hb0ca: y = 16'hfe00;
			16'hb0cb: y = 16'hfe00;
			16'hb0cc: y = 16'hfe00;
			16'hb0cd: y = 16'hfe00;
			16'hb0ce: y = 16'hfe00;
			16'hb0cf: y = 16'hfe00;
			16'hb0d0: y = 16'hfe00;
			16'hb0d1: y = 16'hfe00;
			16'hb0d2: y = 16'hfe00;
			16'hb0d3: y = 16'hfe00;
			16'hb0d4: y = 16'hfe00;
			16'hb0d5: y = 16'hfe00;
			16'hb0d6: y = 16'hfe00;
			16'hb0d7: y = 16'hfe00;
			16'hb0d8: y = 16'hfe00;
			16'hb0d9: y = 16'hfe00;
			16'hb0da: y = 16'hfe00;
			16'hb0db: y = 16'hfe00;
			16'hb0dc: y = 16'hfe00;
			16'hb0dd: y = 16'hfe00;
			16'hb0de: y = 16'hfe00;
			16'hb0df: y = 16'hfe00;
			16'hb0e0: y = 16'hfe00;
			16'hb0e1: y = 16'hfe00;
			16'hb0e2: y = 16'hfe00;
			16'hb0e3: y = 16'hfe00;
			16'hb0e4: y = 16'hfe00;
			16'hb0e5: y = 16'hfe00;
			16'hb0e6: y = 16'hfe00;
			16'hb0e7: y = 16'hfe00;
			16'hb0e8: y = 16'hfe00;
			16'hb0e9: y = 16'hfe00;
			16'hb0ea: y = 16'hfe00;
			16'hb0eb: y = 16'hfe00;
			16'hb0ec: y = 16'hfe00;
			16'hb0ed: y = 16'hfe00;
			16'hb0ee: y = 16'hfe00;
			16'hb0ef: y = 16'hfe00;
			16'hb0f0: y = 16'hfe00;
			16'hb0f1: y = 16'hfe00;
			16'hb0f2: y = 16'hfe00;
			16'hb0f3: y = 16'hfe00;
			16'hb0f4: y = 16'hfe00;
			16'hb0f5: y = 16'hfe00;
			16'hb0f6: y = 16'hfe00;
			16'hb0f7: y = 16'hfe00;
			16'hb0f8: y = 16'hfe00;
			16'hb0f9: y = 16'hfe00;
			16'hb0fa: y = 16'hfe00;
			16'hb0fb: y = 16'hfe00;
			16'hb0fc: y = 16'hfe00;
			16'hb0fd: y = 16'hfe00;
			16'hb0fe: y = 16'hfe00;
			16'hb0ff: y = 16'hfe00;
			16'hb100: y = 16'hfe00;
			16'hb101: y = 16'hfe00;
			16'hb102: y = 16'hfe00;
			16'hb103: y = 16'hfe00;
			16'hb104: y = 16'hfe00;
			16'hb105: y = 16'hfe00;
			16'hb106: y = 16'hfe00;
			16'hb107: y = 16'hfe00;
			16'hb108: y = 16'hfe00;
			16'hb109: y = 16'hfe00;
			16'hb10a: y = 16'hfe00;
			16'hb10b: y = 16'hfe00;
			16'hb10c: y = 16'hfe00;
			16'hb10d: y = 16'hfe00;
			16'hb10e: y = 16'hfe00;
			16'hb10f: y = 16'hfe00;
			16'hb110: y = 16'hfe00;
			16'hb111: y = 16'hfe00;
			16'hb112: y = 16'hfe00;
			16'hb113: y = 16'hfe00;
			16'hb114: y = 16'hfe00;
			16'hb115: y = 16'hfe00;
			16'hb116: y = 16'hfe00;
			16'hb117: y = 16'hfe00;
			16'hb118: y = 16'hfe00;
			16'hb119: y = 16'hfe00;
			16'hb11a: y = 16'hfe00;
			16'hb11b: y = 16'hfe00;
			16'hb11c: y = 16'hfe00;
			16'hb11d: y = 16'hfe00;
			16'hb11e: y = 16'hfe00;
			16'hb11f: y = 16'hfe00;
			16'hb120: y = 16'hfe00;
			16'hb121: y = 16'hfe00;
			16'hb122: y = 16'hfe00;
			16'hb123: y = 16'hfe00;
			16'hb124: y = 16'hfe00;
			16'hb125: y = 16'hfe00;
			16'hb126: y = 16'hfe00;
			16'hb127: y = 16'hfe00;
			16'hb128: y = 16'hfe00;
			16'hb129: y = 16'hfe00;
			16'hb12a: y = 16'hfe00;
			16'hb12b: y = 16'hfe00;
			16'hb12c: y = 16'hfe00;
			16'hb12d: y = 16'hfe00;
			16'hb12e: y = 16'hfe00;
			16'hb12f: y = 16'hfe00;
			16'hb130: y = 16'hfe00;
			16'hb131: y = 16'hfe00;
			16'hb132: y = 16'hfe00;
			16'hb133: y = 16'hfe00;
			16'hb134: y = 16'hfe00;
			16'hb135: y = 16'hfe00;
			16'hb136: y = 16'hfe00;
			16'hb137: y = 16'hfe00;
			16'hb138: y = 16'hfe00;
			16'hb139: y = 16'hfe00;
			16'hb13a: y = 16'hfe00;
			16'hb13b: y = 16'hfe00;
			16'hb13c: y = 16'hfe00;
			16'hb13d: y = 16'hfe00;
			16'hb13e: y = 16'hfe00;
			16'hb13f: y = 16'hfe00;
			16'hb140: y = 16'hfe00;
			16'hb141: y = 16'hfe00;
			16'hb142: y = 16'hfe00;
			16'hb143: y = 16'hfe00;
			16'hb144: y = 16'hfe00;
			16'hb145: y = 16'hfe00;
			16'hb146: y = 16'hfe00;
			16'hb147: y = 16'hfe00;
			16'hb148: y = 16'hfe00;
			16'hb149: y = 16'hfe00;
			16'hb14a: y = 16'hfe00;
			16'hb14b: y = 16'hfe00;
			16'hb14c: y = 16'hfe00;
			16'hb14d: y = 16'hfe00;
			16'hb14e: y = 16'hfe00;
			16'hb14f: y = 16'hfe00;
			16'hb150: y = 16'hfe00;
			16'hb151: y = 16'hfe00;
			16'hb152: y = 16'hfe00;
			16'hb153: y = 16'hfe00;
			16'hb154: y = 16'hfe00;
			16'hb155: y = 16'hfe00;
			16'hb156: y = 16'hfe00;
			16'hb157: y = 16'hfe00;
			16'hb158: y = 16'hfe00;
			16'hb159: y = 16'hfe00;
			16'hb15a: y = 16'hfe00;
			16'hb15b: y = 16'hfe00;
			16'hb15c: y = 16'hfe00;
			16'hb15d: y = 16'hfe00;
			16'hb15e: y = 16'hfe00;
			16'hb15f: y = 16'hfe00;
			16'hb160: y = 16'hfe00;
			16'hb161: y = 16'hfe00;
			16'hb162: y = 16'hfe00;
			16'hb163: y = 16'hfe00;
			16'hb164: y = 16'hfe00;
			16'hb165: y = 16'hfe00;
			16'hb166: y = 16'hfe00;
			16'hb167: y = 16'hfe00;
			16'hb168: y = 16'hfe00;
			16'hb169: y = 16'hfe00;
			16'hb16a: y = 16'hfe00;
			16'hb16b: y = 16'hfe00;
			16'hb16c: y = 16'hfe00;
			16'hb16d: y = 16'hfe00;
			16'hb16e: y = 16'hfe00;
			16'hb16f: y = 16'hfe00;
			16'hb170: y = 16'hfe00;
			16'hb171: y = 16'hfe00;
			16'hb172: y = 16'hfe00;
			16'hb173: y = 16'hfe00;
			16'hb174: y = 16'hfe00;
			16'hb175: y = 16'hfe00;
			16'hb176: y = 16'hfe00;
			16'hb177: y = 16'hfe00;
			16'hb178: y = 16'hfe00;
			16'hb179: y = 16'hfe00;
			16'hb17a: y = 16'hfe00;
			16'hb17b: y = 16'hfe00;
			16'hb17c: y = 16'hfe00;
			16'hb17d: y = 16'hfe00;
			16'hb17e: y = 16'hfe00;
			16'hb17f: y = 16'hfe00;
			16'hb180: y = 16'hfe00;
			16'hb181: y = 16'hfe00;
			16'hb182: y = 16'hfe00;
			16'hb183: y = 16'hfe00;
			16'hb184: y = 16'hfe00;
			16'hb185: y = 16'hfe00;
			16'hb186: y = 16'hfe00;
			16'hb187: y = 16'hfe00;
			16'hb188: y = 16'hfe00;
			16'hb189: y = 16'hfe00;
			16'hb18a: y = 16'hfe00;
			16'hb18b: y = 16'hfe00;
			16'hb18c: y = 16'hfe00;
			16'hb18d: y = 16'hfe00;
			16'hb18e: y = 16'hfe00;
			16'hb18f: y = 16'hfe00;
			16'hb190: y = 16'hfe00;
			16'hb191: y = 16'hfe00;
			16'hb192: y = 16'hfe00;
			16'hb193: y = 16'hfe00;
			16'hb194: y = 16'hfe00;
			16'hb195: y = 16'hfe00;
			16'hb196: y = 16'hfe00;
			16'hb197: y = 16'hfe00;
			16'hb198: y = 16'hfe00;
			16'hb199: y = 16'hfe00;
			16'hb19a: y = 16'hfe00;
			16'hb19b: y = 16'hfe00;
			16'hb19c: y = 16'hfe00;
			16'hb19d: y = 16'hfe00;
			16'hb19e: y = 16'hfe00;
			16'hb19f: y = 16'hfe00;
			16'hb1a0: y = 16'hfe00;
			16'hb1a1: y = 16'hfe00;
			16'hb1a2: y = 16'hfe00;
			16'hb1a3: y = 16'hfe00;
			16'hb1a4: y = 16'hfe00;
			16'hb1a5: y = 16'hfe00;
			16'hb1a6: y = 16'hfe00;
			16'hb1a7: y = 16'hfe00;
			16'hb1a8: y = 16'hfe00;
			16'hb1a9: y = 16'hfe00;
			16'hb1aa: y = 16'hfe00;
			16'hb1ab: y = 16'hfe00;
			16'hb1ac: y = 16'hfe00;
			16'hb1ad: y = 16'hfe00;
			16'hb1ae: y = 16'hfe00;
			16'hb1af: y = 16'hfe00;
			16'hb1b0: y = 16'hfe00;
			16'hb1b1: y = 16'hfe00;
			16'hb1b2: y = 16'hfe00;
			16'hb1b3: y = 16'hfe00;
			16'hb1b4: y = 16'hfe00;
			16'hb1b5: y = 16'hfe00;
			16'hb1b6: y = 16'hfe00;
			16'hb1b7: y = 16'hfe00;
			16'hb1b8: y = 16'hfe00;
			16'hb1b9: y = 16'hfe00;
			16'hb1ba: y = 16'hfe00;
			16'hb1bb: y = 16'hfe00;
			16'hb1bc: y = 16'hfe00;
			16'hb1bd: y = 16'hfe00;
			16'hb1be: y = 16'hfe00;
			16'hb1bf: y = 16'hfe00;
			16'hb1c0: y = 16'hfe00;
			16'hb1c1: y = 16'hfe00;
			16'hb1c2: y = 16'hfe00;
			16'hb1c3: y = 16'hfe00;
			16'hb1c4: y = 16'hfe00;
			16'hb1c5: y = 16'hfe00;
			16'hb1c6: y = 16'hfe00;
			16'hb1c7: y = 16'hfe00;
			16'hb1c8: y = 16'hfe00;
			16'hb1c9: y = 16'hfe00;
			16'hb1ca: y = 16'hfe00;
			16'hb1cb: y = 16'hfe00;
			16'hb1cc: y = 16'hfe00;
			16'hb1cd: y = 16'hfe00;
			16'hb1ce: y = 16'hfe00;
			16'hb1cf: y = 16'hfe00;
			16'hb1d0: y = 16'hfe00;
			16'hb1d1: y = 16'hfe00;
			16'hb1d2: y = 16'hfe00;
			16'hb1d3: y = 16'hfe00;
			16'hb1d4: y = 16'hfe00;
			16'hb1d5: y = 16'hfe00;
			16'hb1d6: y = 16'hfe00;
			16'hb1d7: y = 16'hfe00;
			16'hb1d8: y = 16'hfe00;
			16'hb1d9: y = 16'hfe00;
			16'hb1da: y = 16'hfe00;
			16'hb1db: y = 16'hfe00;
			16'hb1dc: y = 16'hfe00;
			16'hb1dd: y = 16'hfe00;
			16'hb1de: y = 16'hfe00;
			16'hb1df: y = 16'hfe00;
			16'hb1e0: y = 16'hfe00;
			16'hb1e1: y = 16'hfe00;
			16'hb1e2: y = 16'hfe00;
			16'hb1e3: y = 16'hfe00;
			16'hb1e4: y = 16'hfe00;
			16'hb1e5: y = 16'hfe00;
			16'hb1e6: y = 16'hfe00;
			16'hb1e7: y = 16'hfe00;
			16'hb1e8: y = 16'hfe00;
			16'hb1e9: y = 16'hfe00;
			16'hb1ea: y = 16'hfe00;
			16'hb1eb: y = 16'hfe00;
			16'hb1ec: y = 16'hfe00;
			16'hb1ed: y = 16'hfe00;
			16'hb1ee: y = 16'hfe00;
			16'hb1ef: y = 16'hfe00;
			16'hb1f0: y = 16'hfe00;
			16'hb1f1: y = 16'hfe00;
			16'hb1f2: y = 16'hfe00;
			16'hb1f3: y = 16'hfe00;
			16'hb1f4: y = 16'hfe00;
			16'hb1f5: y = 16'hfe00;
			16'hb1f6: y = 16'hfe00;
			16'hb1f7: y = 16'hfe00;
			16'hb1f8: y = 16'hfe00;
			16'hb1f9: y = 16'hfe00;
			16'hb1fa: y = 16'hfe00;
			16'hb1fb: y = 16'hfe00;
			16'hb1fc: y = 16'hfe00;
			16'hb1fd: y = 16'hfe00;
			16'hb1fe: y = 16'hfe00;
			16'hb1ff: y = 16'hfe00;
			16'hb200: y = 16'hfe00;
			16'hb201: y = 16'hfe00;
			16'hb202: y = 16'hfe00;
			16'hb203: y = 16'hfe00;
			16'hb204: y = 16'hfe00;
			16'hb205: y = 16'hfe00;
			16'hb206: y = 16'hfe00;
			16'hb207: y = 16'hfe00;
			16'hb208: y = 16'hfe00;
			16'hb209: y = 16'hfe00;
			16'hb20a: y = 16'hfe00;
			16'hb20b: y = 16'hfe00;
			16'hb20c: y = 16'hfe00;
			16'hb20d: y = 16'hfe00;
			16'hb20e: y = 16'hfe00;
			16'hb20f: y = 16'hfe00;
			16'hb210: y = 16'hfe00;
			16'hb211: y = 16'hfe00;
			16'hb212: y = 16'hfe00;
			16'hb213: y = 16'hfe00;
			16'hb214: y = 16'hfe00;
			16'hb215: y = 16'hfe00;
			16'hb216: y = 16'hfe00;
			16'hb217: y = 16'hfe00;
			16'hb218: y = 16'hfe00;
			16'hb219: y = 16'hfe00;
			16'hb21a: y = 16'hfe00;
			16'hb21b: y = 16'hfe00;
			16'hb21c: y = 16'hfe00;
			16'hb21d: y = 16'hfe00;
			16'hb21e: y = 16'hfe00;
			16'hb21f: y = 16'hfe00;
			16'hb220: y = 16'hfe00;
			16'hb221: y = 16'hfe00;
			16'hb222: y = 16'hfe00;
			16'hb223: y = 16'hfe00;
			16'hb224: y = 16'hfe00;
			16'hb225: y = 16'hfe00;
			16'hb226: y = 16'hfe00;
			16'hb227: y = 16'hfe00;
			16'hb228: y = 16'hfe00;
			16'hb229: y = 16'hfe00;
			16'hb22a: y = 16'hfe00;
			16'hb22b: y = 16'hfe00;
			16'hb22c: y = 16'hfe00;
			16'hb22d: y = 16'hfe00;
			16'hb22e: y = 16'hfe00;
			16'hb22f: y = 16'hfe00;
			16'hb230: y = 16'hfe00;
			16'hb231: y = 16'hfe00;
			16'hb232: y = 16'hfe00;
			16'hb233: y = 16'hfe00;
			16'hb234: y = 16'hfe00;
			16'hb235: y = 16'hfe00;
			16'hb236: y = 16'hfe00;
			16'hb237: y = 16'hfe00;
			16'hb238: y = 16'hfe00;
			16'hb239: y = 16'hfe00;
			16'hb23a: y = 16'hfe00;
			16'hb23b: y = 16'hfe00;
			16'hb23c: y = 16'hfe00;
			16'hb23d: y = 16'hfe00;
			16'hb23e: y = 16'hfe00;
			16'hb23f: y = 16'hfe00;
			16'hb240: y = 16'hfe00;
			16'hb241: y = 16'hfe00;
			16'hb242: y = 16'hfe00;
			16'hb243: y = 16'hfe00;
			16'hb244: y = 16'hfe00;
			16'hb245: y = 16'hfe00;
			16'hb246: y = 16'hfe00;
			16'hb247: y = 16'hfe00;
			16'hb248: y = 16'hfe00;
			16'hb249: y = 16'hfe00;
			16'hb24a: y = 16'hfe00;
			16'hb24b: y = 16'hfe00;
			16'hb24c: y = 16'hfe00;
			16'hb24d: y = 16'hfe00;
			16'hb24e: y = 16'hfe00;
			16'hb24f: y = 16'hfe00;
			16'hb250: y = 16'hfe00;
			16'hb251: y = 16'hfe00;
			16'hb252: y = 16'hfe00;
			16'hb253: y = 16'hfe00;
			16'hb254: y = 16'hfe00;
			16'hb255: y = 16'hfe00;
			16'hb256: y = 16'hfe00;
			16'hb257: y = 16'hfe00;
			16'hb258: y = 16'hfe00;
			16'hb259: y = 16'hfe00;
			16'hb25a: y = 16'hfe00;
			16'hb25b: y = 16'hfe00;
			16'hb25c: y = 16'hfe00;
			16'hb25d: y = 16'hfe00;
			16'hb25e: y = 16'hfe00;
			16'hb25f: y = 16'hfe00;
			16'hb260: y = 16'hfe00;
			16'hb261: y = 16'hfe00;
			16'hb262: y = 16'hfe00;
			16'hb263: y = 16'hfe00;
			16'hb264: y = 16'hfe00;
			16'hb265: y = 16'hfe00;
			16'hb266: y = 16'hfe00;
			16'hb267: y = 16'hfe00;
			16'hb268: y = 16'hfe00;
			16'hb269: y = 16'hfe00;
			16'hb26a: y = 16'hfe00;
			16'hb26b: y = 16'hfe00;
			16'hb26c: y = 16'hfe00;
			16'hb26d: y = 16'hfe00;
			16'hb26e: y = 16'hfe00;
			16'hb26f: y = 16'hfe00;
			16'hb270: y = 16'hfe00;
			16'hb271: y = 16'hfe00;
			16'hb272: y = 16'hfe00;
			16'hb273: y = 16'hfe00;
			16'hb274: y = 16'hfe00;
			16'hb275: y = 16'hfe00;
			16'hb276: y = 16'hfe00;
			16'hb277: y = 16'hfe00;
			16'hb278: y = 16'hfe00;
			16'hb279: y = 16'hfe00;
			16'hb27a: y = 16'hfe00;
			16'hb27b: y = 16'hfe00;
			16'hb27c: y = 16'hfe00;
			16'hb27d: y = 16'hfe00;
			16'hb27e: y = 16'hfe00;
			16'hb27f: y = 16'hfe00;
			16'hb280: y = 16'hfe00;
			16'hb281: y = 16'hfe00;
			16'hb282: y = 16'hfe00;
			16'hb283: y = 16'hfe00;
			16'hb284: y = 16'hfe00;
			16'hb285: y = 16'hfe00;
			16'hb286: y = 16'hfe00;
			16'hb287: y = 16'hfe00;
			16'hb288: y = 16'hfe00;
			16'hb289: y = 16'hfe00;
			16'hb28a: y = 16'hfe00;
			16'hb28b: y = 16'hfe00;
			16'hb28c: y = 16'hfe00;
			16'hb28d: y = 16'hfe00;
			16'hb28e: y = 16'hfe00;
			16'hb28f: y = 16'hfe00;
			16'hb290: y = 16'hfe00;
			16'hb291: y = 16'hfe00;
			16'hb292: y = 16'hfe00;
			16'hb293: y = 16'hfe00;
			16'hb294: y = 16'hfe00;
			16'hb295: y = 16'hfe00;
			16'hb296: y = 16'hfe00;
			16'hb297: y = 16'hfe00;
			16'hb298: y = 16'hfe00;
			16'hb299: y = 16'hfe00;
			16'hb29a: y = 16'hfe00;
			16'hb29b: y = 16'hfe00;
			16'hb29c: y = 16'hfe00;
			16'hb29d: y = 16'hfe00;
			16'hb29e: y = 16'hfe00;
			16'hb29f: y = 16'hfe00;
			16'hb2a0: y = 16'hfe00;
			16'hb2a1: y = 16'hfe00;
			16'hb2a2: y = 16'hfe00;
			16'hb2a3: y = 16'hfe00;
			16'hb2a4: y = 16'hfe00;
			16'hb2a5: y = 16'hfe00;
			16'hb2a6: y = 16'hfe00;
			16'hb2a7: y = 16'hfe00;
			16'hb2a8: y = 16'hfe00;
			16'hb2a9: y = 16'hfe00;
			16'hb2aa: y = 16'hfe00;
			16'hb2ab: y = 16'hfe00;
			16'hb2ac: y = 16'hfe00;
			16'hb2ad: y = 16'hfe00;
			16'hb2ae: y = 16'hfe00;
			16'hb2af: y = 16'hfe00;
			16'hb2b0: y = 16'hfe00;
			16'hb2b1: y = 16'hfe00;
			16'hb2b2: y = 16'hfe00;
			16'hb2b3: y = 16'hfe00;
			16'hb2b4: y = 16'hfe00;
			16'hb2b5: y = 16'hfe00;
			16'hb2b6: y = 16'hfe00;
			16'hb2b7: y = 16'hfe00;
			16'hb2b8: y = 16'hfe00;
			16'hb2b9: y = 16'hfe00;
			16'hb2ba: y = 16'hfe00;
			16'hb2bb: y = 16'hfe00;
			16'hb2bc: y = 16'hfe00;
			16'hb2bd: y = 16'hfe00;
			16'hb2be: y = 16'hfe00;
			16'hb2bf: y = 16'hfe00;
			16'hb2c0: y = 16'hfe00;
			16'hb2c1: y = 16'hfe00;
			16'hb2c2: y = 16'hfe00;
			16'hb2c3: y = 16'hfe00;
			16'hb2c4: y = 16'hfe00;
			16'hb2c5: y = 16'hfe00;
			16'hb2c6: y = 16'hfe00;
			16'hb2c7: y = 16'hfe00;
			16'hb2c8: y = 16'hfe00;
			16'hb2c9: y = 16'hfe00;
			16'hb2ca: y = 16'hfe00;
			16'hb2cb: y = 16'hfe00;
			16'hb2cc: y = 16'hfe00;
			16'hb2cd: y = 16'hfe00;
			16'hb2ce: y = 16'hfe00;
			16'hb2cf: y = 16'hfe00;
			16'hb2d0: y = 16'hfe00;
			16'hb2d1: y = 16'hfe00;
			16'hb2d2: y = 16'hfe00;
			16'hb2d3: y = 16'hfe00;
			16'hb2d4: y = 16'hfe00;
			16'hb2d5: y = 16'hfe00;
			16'hb2d6: y = 16'hfe00;
			16'hb2d7: y = 16'hfe00;
			16'hb2d8: y = 16'hfe00;
			16'hb2d9: y = 16'hfe00;
			16'hb2da: y = 16'hfe00;
			16'hb2db: y = 16'hfe00;
			16'hb2dc: y = 16'hfe00;
			16'hb2dd: y = 16'hfe00;
			16'hb2de: y = 16'hfe00;
			16'hb2df: y = 16'hfe00;
			16'hb2e0: y = 16'hfe00;
			16'hb2e1: y = 16'hfe00;
			16'hb2e2: y = 16'hfe00;
			16'hb2e3: y = 16'hfe00;
			16'hb2e4: y = 16'hfe00;
			16'hb2e5: y = 16'hfe00;
			16'hb2e6: y = 16'hfe00;
			16'hb2e7: y = 16'hfe00;
			16'hb2e8: y = 16'hfe00;
			16'hb2e9: y = 16'hfe00;
			16'hb2ea: y = 16'hfe00;
			16'hb2eb: y = 16'hfe00;
			16'hb2ec: y = 16'hfe00;
			16'hb2ed: y = 16'hfe00;
			16'hb2ee: y = 16'hfe00;
			16'hb2ef: y = 16'hfe00;
			16'hb2f0: y = 16'hfe00;
			16'hb2f1: y = 16'hfe00;
			16'hb2f2: y = 16'hfe00;
			16'hb2f3: y = 16'hfe00;
			16'hb2f4: y = 16'hfe00;
			16'hb2f5: y = 16'hfe00;
			16'hb2f6: y = 16'hfe00;
			16'hb2f7: y = 16'hfe00;
			16'hb2f8: y = 16'hfe00;
			16'hb2f9: y = 16'hfe00;
			16'hb2fa: y = 16'hfe00;
			16'hb2fb: y = 16'hfe00;
			16'hb2fc: y = 16'hfe00;
			16'hb2fd: y = 16'hfe00;
			16'hb2fe: y = 16'hfe00;
			16'hb2ff: y = 16'hfe00;
			16'hb300: y = 16'hfe00;
			16'hb301: y = 16'hfe00;
			16'hb302: y = 16'hfe00;
			16'hb303: y = 16'hfe00;
			16'hb304: y = 16'hfe00;
			16'hb305: y = 16'hfe00;
			16'hb306: y = 16'hfe00;
			16'hb307: y = 16'hfe00;
			16'hb308: y = 16'hfe00;
			16'hb309: y = 16'hfe00;
			16'hb30a: y = 16'hfe00;
			16'hb30b: y = 16'hfe00;
			16'hb30c: y = 16'hfe00;
			16'hb30d: y = 16'hfe00;
			16'hb30e: y = 16'hfe00;
			16'hb30f: y = 16'hfe00;
			16'hb310: y = 16'hfe00;
			16'hb311: y = 16'hfe00;
			16'hb312: y = 16'hfe00;
			16'hb313: y = 16'hfe00;
			16'hb314: y = 16'hfe00;
			16'hb315: y = 16'hfe00;
			16'hb316: y = 16'hfe00;
			16'hb317: y = 16'hfe00;
			16'hb318: y = 16'hfe00;
			16'hb319: y = 16'hfe00;
			16'hb31a: y = 16'hfe00;
			16'hb31b: y = 16'hfe00;
			16'hb31c: y = 16'hfe00;
			16'hb31d: y = 16'hfe00;
			16'hb31e: y = 16'hfe00;
			16'hb31f: y = 16'hfe00;
			16'hb320: y = 16'hfe00;
			16'hb321: y = 16'hfe00;
			16'hb322: y = 16'hfe00;
			16'hb323: y = 16'hfe00;
			16'hb324: y = 16'hfe00;
			16'hb325: y = 16'hfe00;
			16'hb326: y = 16'hfe00;
			16'hb327: y = 16'hfe00;
			16'hb328: y = 16'hfe00;
			16'hb329: y = 16'hfe00;
			16'hb32a: y = 16'hfe00;
			16'hb32b: y = 16'hfe00;
			16'hb32c: y = 16'hfe00;
			16'hb32d: y = 16'hfe00;
			16'hb32e: y = 16'hfe00;
			16'hb32f: y = 16'hfe00;
			16'hb330: y = 16'hfe00;
			16'hb331: y = 16'hfe00;
			16'hb332: y = 16'hfe00;
			16'hb333: y = 16'hfe00;
			16'hb334: y = 16'hfe00;
			16'hb335: y = 16'hfe00;
			16'hb336: y = 16'hfe00;
			16'hb337: y = 16'hfe00;
			16'hb338: y = 16'hfe00;
			16'hb339: y = 16'hfe00;
			16'hb33a: y = 16'hfe00;
			16'hb33b: y = 16'hfe00;
			16'hb33c: y = 16'hfe00;
			16'hb33d: y = 16'hfe00;
			16'hb33e: y = 16'hfe00;
			16'hb33f: y = 16'hfe00;
			16'hb340: y = 16'hfe00;
			16'hb341: y = 16'hfe00;
			16'hb342: y = 16'hfe00;
			16'hb343: y = 16'hfe00;
			16'hb344: y = 16'hfe00;
			16'hb345: y = 16'hfe00;
			16'hb346: y = 16'hfe00;
			16'hb347: y = 16'hfe00;
			16'hb348: y = 16'hfe00;
			16'hb349: y = 16'hfe00;
			16'hb34a: y = 16'hfe00;
			16'hb34b: y = 16'hfe00;
			16'hb34c: y = 16'hfe00;
			16'hb34d: y = 16'hfe00;
			16'hb34e: y = 16'hfe00;
			16'hb34f: y = 16'hfe00;
			16'hb350: y = 16'hfe00;
			16'hb351: y = 16'hfe00;
			16'hb352: y = 16'hfe00;
			16'hb353: y = 16'hfe00;
			16'hb354: y = 16'hfe00;
			16'hb355: y = 16'hfe00;
			16'hb356: y = 16'hfe00;
			16'hb357: y = 16'hfe00;
			16'hb358: y = 16'hfe00;
			16'hb359: y = 16'hfe00;
			16'hb35a: y = 16'hfe00;
			16'hb35b: y = 16'hfe00;
			16'hb35c: y = 16'hfe00;
			16'hb35d: y = 16'hfe00;
			16'hb35e: y = 16'hfe00;
			16'hb35f: y = 16'hfe00;
			16'hb360: y = 16'hfe00;
			16'hb361: y = 16'hfe00;
			16'hb362: y = 16'hfe00;
			16'hb363: y = 16'hfe00;
			16'hb364: y = 16'hfe00;
			16'hb365: y = 16'hfe00;
			16'hb366: y = 16'hfe00;
			16'hb367: y = 16'hfe00;
			16'hb368: y = 16'hfe00;
			16'hb369: y = 16'hfe00;
			16'hb36a: y = 16'hfe00;
			16'hb36b: y = 16'hfe00;
			16'hb36c: y = 16'hfe00;
			16'hb36d: y = 16'hfe00;
			16'hb36e: y = 16'hfe00;
			16'hb36f: y = 16'hfe00;
			16'hb370: y = 16'hfe00;
			16'hb371: y = 16'hfe00;
			16'hb372: y = 16'hfe00;
			16'hb373: y = 16'hfe00;
			16'hb374: y = 16'hfe00;
			16'hb375: y = 16'hfe00;
			16'hb376: y = 16'hfe00;
			16'hb377: y = 16'hfe00;
			16'hb378: y = 16'hfe00;
			16'hb379: y = 16'hfe00;
			16'hb37a: y = 16'hfe00;
			16'hb37b: y = 16'hfe00;
			16'hb37c: y = 16'hfe00;
			16'hb37d: y = 16'hfe00;
			16'hb37e: y = 16'hfe00;
			16'hb37f: y = 16'hfe00;
			16'hb380: y = 16'hfe00;
			16'hb381: y = 16'hfe00;
			16'hb382: y = 16'hfe00;
			16'hb383: y = 16'hfe00;
			16'hb384: y = 16'hfe00;
			16'hb385: y = 16'hfe00;
			16'hb386: y = 16'hfe00;
			16'hb387: y = 16'hfe00;
			16'hb388: y = 16'hfe00;
			16'hb389: y = 16'hfe00;
			16'hb38a: y = 16'hfe00;
			16'hb38b: y = 16'hfe00;
			16'hb38c: y = 16'hfe00;
			16'hb38d: y = 16'hfe00;
			16'hb38e: y = 16'hfe00;
			16'hb38f: y = 16'hfe00;
			16'hb390: y = 16'hfe00;
			16'hb391: y = 16'hfe00;
			16'hb392: y = 16'hfe00;
			16'hb393: y = 16'hfe00;
			16'hb394: y = 16'hfe00;
			16'hb395: y = 16'hfe00;
			16'hb396: y = 16'hfe00;
			16'hb397: y = 16'hfe00;
			16'hb398: y = 16'hfe00;
			16'hb399: y = 16'hfe00;
			16'hb39a: y = 16'hfe00;
			16'hb39b: y = 16'hfe00;
			16'hb39c: y = 16'hfe00;
			16'hb39d: y = 16'hfe00;
			16'hb39e: y = 16'hfe00;
			16'hb39f: y = 16'hfe00;
			16'hb3a0: y = 16'hfe00;
			16'hb3a1: y = 16'hfe00;
			16'hb3a2: y = 16'hfe00;
			16'hb3a3: y = 16'hfe00;
			16'hb3a4: y = 16'hfe00;
			16'hb3a5: y = 16'hfe00;
			16'hb3a6: y = 16'hfe00;
			16'hb3a7: y = 16'hfe00;
			16'hb3a8: y = 16'hfe00;
			16'hb3a9: y = 16'hfe00;
			16'hb3aa: y = 16'hfe00;
			16'hb3ab: y = 16'hfe00;
			16'hb3ac: y = 16'hfe00;
			16'hb3ad: y = 16'hfe00;
			16'hb3ae: y = 16'hfe00;
			16'hb3af: y = 16'hfe00;
			16'hb3b0: y = 16'hfe00;
			16'hb3b1: y = 16'hfe00;
			16'hb3b2: y = 16'hfe00;
			16'hb3b3: y = 16'hfe00;
			16'hb3b4: y = 16'hfe00;
			16'hb3b5: y = 16'hfe00;
			16'hb3b6: y = 16'hfe00;
			16'hb3b7: y = 16'hfe00;
			16'hb3b8: y = 16'hfe00;
			16'hb3b9: y = 16'hfe00;
			16'hb3ba: y = 16'hfe00;
			16'hb3bb: y = 16'hfe00;
			16'hb3bc: y = 16'hfe00;
			16'hb3bd: y = 16'hfe00;
			16'hb3be: y = 16'hfe00;
			16'hb3bf: y = 16'hfe00;
			16'hb3c0: y = 16'hfe00;
			16'hb3c1: y = 16'hfe00;
			16'hb3c2: y = 16'hfe00;
			16'hb3c3: y = 16'hfe00;
			16'hb3c4: y = 16'hfe00;
			16'hb3c5: y = 16'hfe00;
			16'hb3c6: y = 16'hfe00;
			16'hb3c7: y = 16'hfe00;
			16'hb3c8: y = 16'hfe00;
			16'hb3c9: y = 16'hfe00;
			16'hb3ca: y = 16'hfe00;
			16'hb3cb: y = 16'hfe00;
			16'hb3cc: y = 16'hfe00;
			16'hb3cd: y = 16'hfe00;
			16'hb3ce: y = 16'hfe00;
			16'hb3cf: y = 16'hfe00;
			16'hb3d0: y = 16'hfe00;
			16'hb3d1: y = 16'hfe00;
			16'hb3d2: y = 16'hfe00;
			16'hb3d3: y = 16'hfe00;
			16'hb3d4: y = 16'hfe00;
			16'hb3d5: y = 16'hfe00;
			16'hb3d6: y = 16'hfe00;
			16'hb3d7: y = 16'hfe00;
			16'hb3d8: y = 16'hfe00;
			16'hb3d9: y = 16'hfe00;
			16'hb3da: y = 16'hfe00;
			16'hb3db: y = 16'hfe00;
			16'hb3dc: y = 16'hfe00;
			16'hb3dd: y = 16'hfe00;
			16'hb3de: y = 16'hfe00;
			16'hb3df: y = 16'hfe00;
			16'hb3e0: y = 16'hfe00;
			16'hb3e1: y = 16'hfe00;
			16'hb3e2: y = 16'hfe00;
			16'hb3e3: y = 16'hfe00;
			16'hb3e4: y = 16'hfe00;
			16'hb3e5: y = 16'hfe00;
			16'hb3e6: y = 16'hfe00;
			16'hb3e7: y = 16'hfe00;
			16'hb3e8: y = 16'hfe00;
			16'hb3e9: y = 16'hfe00;
			16'hb3ea: y = 16'hfe00;
			16'hb3eb: y = 16'hfe00;
			16'hb3ec: y = 16'hfe00;
			16'hb3ed: y = 16'hfe00;
			16'hb3ee: y = 16'hfe00;
			16'hb3ef: y = 16'hfe00;
			16'hb3f0: y = 16'hfe00;
			16'hb3f1: y = 16'hfe00;
			16'hb3f2: y = 16'hfe00;
			16'hb3f3: y = 16'hfe00;
			16'hb3f4: y = 16'hfe00;
			16'hb3f5: y = 16'hfe00;
			16'hb3f6: y = 16'hfe00;
			16'hb3f7: y = 16'hfe00;
			16'hb3f8: y = 16'hfe00;
			16'hb3f9: y = 16'hfe00;
			16'hb3fa: y = 16'hfe00;
			16'hb3fb: y = 16'hfe00;
			16'hb3fc: y = 16'hfe00;
			16'hb3fd: y = 16'hfe00;
			16'hb3fe: y = 16'hfe00;
			16'hb3ff: y = 16'hfe00;
			16'hb400: y = 16'hfe00;
			16'hb401: y = 16'hfe00;
			16'hb402: y = 16'hfe00;
			16'hb403: y = 16'hfe00;
			16'hb404: y = 16'hfe00;
			16'hb405: y = 16'hfe00;
			16'hb406: y = 16'hfe00;
			16'hb407: y = 16'hfe00;
			16'hb408: y = 16'hfe00;
			16'hb409: y = 16'hfe00;
			16'hb40a: y = 16'hfe00;
			16'hb40b: y = 16'hfe00;
			16'hb40c: y = 16'hfe00;
			16'hb40d: y = 16'hfe00;
			16'hb40e: y = 16'hfe00;
			16'hb40f: y = 16'hfe00;
			16'hb410: y = 16'hfe00;
			16'hb411: y = 16'hfe00;
			16'hb412: y = 16'hfe00;
			16'hb413: y = 16'hfe00;
			16'hb414: y = 16'hfe00;
			16'hb415: y = 16'hfe00;
			16'hb416: y = 16'hfe00;
			16'hb417: y = 16'hfe00;
			16'hb418: y = 16'hfe00;
			16'hb419: y = 16'hfe00;
			16'hb41a: y = 16'hfe00;
			16'hb41b: y = 16'hfe00;
			16'hb41c: y = 16'hfe00;
			16'hb41d: y = 16'hfe00;
			16'hb41e: y = 16'hfe00;
			16'hb41f: y = 16'hfe00;
			16'hb420: y = 16'hfe00;
			16'hb421: y = 16'hfe00;
			16'hb422: y = 16'hfe00;
			16'hb423: y = 16'hfe00;
			16'hb424: y = 16'hfe00;
			16'hb425: y = 16'hfe00;
			16'hb426: y = 16'hfe00;
			16'hb427: y = 16'hfe00;
			16'hb428: y = 16'hfe00;
			16'hb429: y = 16'hfe00;
			16'hb42a: y = 16'hfe00;
			16'hb42b: y = 16'hfe00;
			16'hb42c: y = 16'hfe00;
			16'hb42d: y = 16'hfe00;
			16'hb42e: y = 16'hfe00;
			16'hb42f: y = 16'hfe00;
			16'hb430: y = 16'hfe00;
			16'hb431: y = 16'hfe00;
			16'hb432: y = 16'hfe00;
			16'hb433: y = 16'hfe00;
			16'hb434: y = 16'hfe00;
			16'hb435: y = 16'hfe00;
			16'hb436: y = 16'hfe00;
			16'hb437: y = 16'hfe00;
			16'hb438: y = 16'hfe00;
			16'hb439: y = 16'hfe00;
			16'hb43a: y = 16'hfe00;
			16'hb43b: y = 16'hfe00;
			16'hb43c: y = 16'hfe00;
			16'hb43d: y = 16'hfe00;
			16'hb43e: y = 16'hfe00;
			16'hb43f: y = 16'hfe00;
			16'hb440: y = 16'hfe00;
			16'hb441: y = 16'hfe00;
			16'hb442: y = 16'hfe00;
			16'hb443: y = 16'hfe00;
			16'hb444: y = 16'hfe00;
			16'hb445: y = 16'hfe00;
			16'hb446: y = 16'hfe00;
			16'hb447: y = 16'hfe00;
			16'hb448: y = 16'hfe00;
			16'hb449: y = 16'hfe00;
			16'hb44a: y = 16'hfe00;
			16'hb44b: y = 16'hfe00;
			16'hb44c: y = 16'hfe00;
			16'hb44d: y = 16'hfe00;
			16'hb44e: y = 16'hfe00;
			16'hb44f: y = 16'hfe00;
			16'hb450: y = 16'hfe00;
			16'hb451: y = 16'hfe00;
			16'hb452: y = 16'hfe00;
			16'hb453: y = 16'hfe00;
			16'hb454: y = 16'hfe00;
			16'hb455: y = 16'hfe00;
			16'hb456: y = 16'hfe00;
			16'hb457: y = 16'hfe00;
			16'hb458: y = 16'hfe00;
			16'hb459: y = 16'hfe00;
			16'hb45a: y = 16'hfe00;
			16'hb45b: y = 16'hfe00;
			16'hb45c: y = 16'hfe00;
			16'hb45d: y = 16'hfe00;
			16'hb45e: y = 16'hfe00;
			16'hb45f: y = 16'hfe00;
			16'hb460: y = 16'hfe00;
			16'hb461: y = 16'hfe00;
			16'hb462: y = 16'hfe00;
			16'hb463: y = 16'hfe00;
			16'hb464: y = 16'hfe00;
			16'hb465: y = 16'hfe00;
			16'hb466: y = 16'hfe00;
			16'hb467: y = 16'hfe00;
			16'hb468: y = 16'hfe00;
			16'hb469: y = 16'hfe00;
			16'hb46a: y = 16'hfe00;
			16'hb46b: y = 16'hfe00;
			16'hb46c: y = 16'hfe00;
			16'hb46d: y = 16'hfe00;
			16'hb46e: y = 16'hfe00;
			16'hb46f: y = 16'hfe00;
			16'hb470: y = 16'hfe00;
			16'hb471: y = 16'hfe00;
			16'hb472: y = 16'hfe00;
			16'hb473: y = 16'hfe00;
			16'hb474: y = 16'hfe00;
			16'hb475: y = 16'hfe00;
			16'hb476: y = 16'hfe00;
			16'hb477: y = 16'hfe00;
			16'hb478: y = 16'hfe00;
			16'hb479: y = 16'hfe00;
			16'hb47a: y = 16'hfe00;
			16'hb47b: y = 16'hfe00;
			16'hb47c: y = 16'hfe00;
			16'hb47d: y = 16'hfe00;
			16'hb47e: y = 16'hfe00;
			16'hb47f: y = 16'hfe00;
			16'hb480: y = 16'hfe00;
			16'hb481: y = 16'hfe00;
			16'hb482: y = 16'hfe00;
			16'hb483: y = 16'hfe00;
			16'hb484: y = 16'hfe00;
			16'hb485: y = 16'hfe00;
			16'hb486: y = 16'hfe00;
			16'hb487: y = 16'hfe00;
			16'hb488: y = 16'hfe00;
			16'hb489: y = 16'hfe00;
			16'hb48a: y = 16'hfe00;
			16'hb48b: y = 16'hfe00;
			16'hb48c: y = 16'hfe00;
			16'hb48d: y = 16'hfe00;
			16'hb48e: y = 16'hfe00;
			16'hb48f: y = 16'hfe00;
			16'hb490: y = 16'hfe00;
			16'hb491: y = 16'hfe00;
			16'hb492: y = 16'hfe00;
			16'hb493: y = 16'hfe00;
			16'hb494: y = 16'hfe00;
			16'hb495: y = 16'hfe00;
			16'hb496: y = 16'hfe00;
			16'hb497: y = 16'hfe00;
			16'hb498: y = 16'hfe00;
			16'hb499: y = 16'hfe00;
			16'hb49a: y = 16'hfe00;
			16'hb49b: y = 16'hfe00;
			16'hb49c: y = 16'hfe00;
			16'hb49d: y = 16'hfe00;
			16'hb49e: y = 16'hfe00;
			16'hb49f: y = 16'hfe00;
			16'hb4a0: y = 16'hfe00;
			16'hb4a1: y = 16'hfe00;
			16'hb4a2: y = 16'hfe00;
			16'hb4a3: y = 16'hfe00;
			16'hb4a4: y = 16'hfe00;
			16'hb4a5: y = 16'hfe00;
			16'hb4a6: y = 16'hfe00;
			16'hb4a7: y = 16'hfe00;
			16'hb4a8: y = 16'hfe00;
			16'hb4a9: y = 16'hfe00;
			16'hb4aa: y = 16'hfe00;
			16'hb4ab: y = 16'hfe00;
			16'hb4ac: y = 16'hfe00;
			16'hb4ad: y = 16'hfe00;
			16'hb4ae: y = 16'hfe00;
			16'hb4af: y = 16'hfe00;
			16'hb4b0: y = 16'hfe00;
			16'hb4b1: y = 16'hfe00;
			16'hb4b2: y = 16'hfe00;
			16'hb4b3: y = 16'hfe00;
			16'hb4b4: y = 16'hfe00;
			16'hb4b5: y = 16'hfe00;
			16'hb4b6: y = 16'hfe00;
			16'hb4b7: y = 16'hfe00;
			16'hb4b8: y = 16'hfe00;
			16'hb4b9: y = 16'hfe00;
			16'hb4ba: y = 16'hfe00;
			16'hb4bb: y = 16'hfe00;
			16'hb4bc: y = 16'hfe00;
			16'hb4bd: y = 16'hfe00;
			16'hb4be: y = 16'hfe00;
			16'hb4bf: y = 16'hfe00;
			16'hb4c0: y = 16'hfe00;
			16'hb4c1: y = 16'hfe00;
			16'hb4c2: y = 16'hfe00;
			16'hb4c3: y = 16'hfe00;
			16'hb4c4: y = 16'hfe00;
			16'hb4c5: y = 16'hfe00;
			16'hb4c6: y = 16'hfe00;
			16'hb4c7: y = 16'hfe00;
			16'hb4c8: y = 16'hfe00;
			16'hb4c9: y = 16'hfe00;
			16'hb4ca: y = 16'hfe00;
			16'hb4cb: y = 16'hfe00;
			16'hb4cc: y = 16'hfe00;
			16'hb4cd: y = 16'hfe00;
			16'hb4ce: y = 16'hfe00;
			16'hb4cf: y = 16'hfe00;
			16'hb4d0: y = 16'hfe00;
			16'hb4d1: y = 16'hfe00;
			16'hb4d2: y = 16'hfe00;
			16'hb4d3: y = 16'hfe00;
			16'hb4d4: y = 16'hfe00;
			16'hb4d5: y = 16'hfe00;
			16'hb4d6: y = 16'hfe00;
			16'hb4d7: y = 16'hfe00;
			16'hb4d8: y = 16'hfe00;
			16'hb4d9: y = 16'hfe00;
			16'hb4da: y = 16'hfe00;
			16'hb4db: y = 16'hfe00;
			16'hb4dc: y = 16'hfe00;
			16'hb4dd: y = 16'hfe00;
			16'hb4de: y = 16'hfe00;
			16'hb4df: y = 16'hfe00;
			16'hb4e0: y = 16'hfe00;
			16'hb4e1: y = 16'hfe00;
			16'hb4e2: y = 16'hfe00;
			16'hb4e3: y = 16'hfe00;
			16'hb4e4: y = 16'hfe00;
			16'hb4e5: y = 16'hfe00;
			16'hb4e6: y = 16'hfe00;
			16'hb4e7: y = 16'hfe00;
			16'hb4e8: y = 16'hfe00;
			16'hb4e9: y = 16'hfe00;
			16'hb4ea: y = 16'hfe00;
			16'hb4eb: y = 16'hfe00;
			16'hb4ec: y = 16'hfe00;
			16'hb4ed: y = 16'hfe00;
			16'hb4ee: y = 16'hfe00;
			16'hb4ef: y = 16'hfe00;
			16'hb4f0: y = 16'hfe00;
			16'hb4f1: y = 16'hfe00;
			16'hb4f2: y = 16'hfe00;
			16'hb4f3: y = 16'hfe00;
			16'hb4f4: y = 16'hfe00;
			16'hb4f5: y = 16'hfe00;
			16'hb4f6: y = 16'hfe00;
			16'hb4f7: y = 16'hfe00;
			16'hb4f8: y = 16'hfe00;
			16'hb4f9: y = 16'hfe00;
			16'hb4fa: y = 16'hfe00;
			16'hb4fb: y = 16'hfe00;
			16'hb4fc: y = 16'hfe00;
			16'hb4fd: y = 16'hfe00;
			16'hb4fe: y = 16'hfe00;
			16'hb4ff: y = 16'hfe00;
			16'hb500: y = 16'hfe00;
			16'hb501: y = 16'hfe00;
			16'hb502: y = 16'hfe00;
			16'hb503: y = 16'hfe00;
			16'hb504: y = 16'hfe00;
			16'hb505: y = 16'hfe00;
			16'hb506: y = 16'hfe00;
			16'hb507: y = 16'hfe00;
			16'hb508: y = 16'hfe00;
			16'hb509: y = 16'hfe00;
			16'hb50a: y = 16'hfe00;
			16'hb50b: y = 16'hfe00;
			16'hb50c: y = 16'hfe00;
			16'hb50d: y = 16'hfe00;
			16'hb50e: y = 16'hfe00;
			16'hb50f: y = 16'hfe00;
			16'hb510: y = 16'hfe00;
			16'hb511: y = 16'hfe00;
			16'hb512: y = 16'hfe00;
			16'hb513: y = 16'hfe00;
			16'hb514: y = 16'hfe00;
			16'hb515: y = 16'hfe00;
			16'hb516: y = 16'hfe00;
			16'hb517: y = 16'hfe00;
			16'hb518: y = 16'hfe00;
			16'hb519: y = 16'hfe00;
			16'hb51a: y = 16'hfe00;
			16'hb51b: y = 16'hfe00;
			16'hb51c: y = 16'hfe00;
			16'hb51d: y = 16'hfe00;
			16'hb51e: y = 16'hfe00;
			16'hb51f: y = 16'hfe00;
			16'hb520: y = 16'hfe00;
			16'hb521: y = 16'hfe00;
			16'hb522: y = 16'hfe00;
			16'hb523: y = 16'hfe00;
			16'hb524: y = 16'hfe00;
			16'hb525: y = 16'hfe00;
			16'hb526: y = 16'hfe00;
			16'hb527: y = 16'hfe00;
			16'hb528: y = 16'hfe00;
			16'hb529: y = 16'hfe00;
			16'hb52a: y = 16'hfe00;
			16'hb52b: y = 16'hfe00;
			16'hb52c: y = 16'hfe00;
			16'hb52d: y = 16'hfe00;
			16'hb52e: y = 16'hfe00;
			16'hb52f: y = 16'hfe00;
			16'hb530: y = 16'hfe00;
			16'hb531: y = 16'hfe00;
			16'hb532: y = 16'hfe00;
			16'hb533: y = 16'hfe00;
			16'hb534: y = 16'hfe00;
			16'hb535: y = 16'hfe00;
			16'hb536: y = 16'hfe00;
			16'hb537: y = 16'hfe00;
			16'hb538: y = 16'hfe00;
			16'hb539: y = 16'hfe00;
			16'hb53a: y = 16'hfe00;
			16'hb53b: y = 16'hfe00;
			16'hb53c: y = 16'hfe00;
			16'hb53d: y = 16'hfe00;
			16'hb53e: y = 16'hfe00;
			16'hb53f: y = 16'hfe00;
			16'hb540: y = 16'hfe00;
			16'hb541: y = 16'hfe00;
			16'hb542: y = 16'hfe00;
			16'hb543: y = 16'hfe00;
			16'hb544: y = 16'hfe00;
			16'hb545: y = 16'hfe00;
			16'hb546: y = 16'hfe00;
			16'hb547: y = 16'hfe00;
			16'hb548: y = 16'hfe00;
			16'hb549: y = 16'hfe00;
			16'hb54a: y = 16'hfe00;
			16'hb54b: y = 16'hfe00;
			16'hb54c: y = 16'hfe00;
			16'hb54d: y = 16'hfe00;
			16'hb54e: y = 16'hfe00;
			16'hb54f: y = 16'hfe00;
			16'hb550: y = 16'hfe00;
			16'hb551: y = 16'hfe00;
			16'hb552: y = 16'hfe00;
			16'hb553: y = 16'hfe00;
			16'hb554: y = 16'hfe00;
			16'hb555: y = 16'hfe00;
			16'hb556: y = 16'hfe00;
			16'hb557: y = 16'hfe00;
			16'hb558: y = 16'hfe00;
			16'hb559: y = 16'hfe00;
			16'hb55a: y = 16'hfe00;
			16'hb55b: y = 16'hfe00;
			16'hb55c: y = 16'hfe00;
			16'hb55d: y = 16'hfe00;
			16'hb55e: y = 16'hfe00;
			16'hb55f: y = 16'hfe00;
			16'hb560: y = 16'hfe00;
			16'hb561: y = 16'hfe00;
			16'hb562: y = 16'hfe00;
			16'hb563: y = 16'hfe00;
			16'hb564: y = 16'hfe00;
			16'hb565: y = 16'hfe00;
			16'hb566: y = 16'hfe00;
			16'hb567: y = 16'hfe00;
			16'hb568: y = 16'hfe00;
			16'hb569: y = 16'hfe00;
			16'hb56a: y = 16'hfe00;
			16'hb56b: y = 16'hfe00;
			16'hb56c: y = 16'hfe00;
			16'hb56d: y = 16'hfe00;
			16'hb56e: y = 16'hfe00;
			16'hb56f: y = 16'hfe00;
			16'hb570: y = 16'hfe00;
			16'hb571: y = 16'hfe00;
			16'hb572: y = 16'hfe00;
			16'hb573: y = 16'hfe00;
			16'hb574: y = 16'hfe00;
			16'hb575: y = 16'hfe00;
			16'hb576: y = 16'hfe00;
			16'hb577: y = 16'hfe00;
			16'hb578: y = 16'hfe00;
			16'hb579: y = 16'hfe00;
			16'hb57a: y = 16'hfe00;
			16'hb57b: y = 16'hfe00;
			16'hb57c: y = 16'hfe00;
			16'hb57d: y = 16'hfe00;
			16'hb57e: y = 16'hfe00;
			16'hb57f: y = 16'hfe00;
			16'hb580: y = 16'hfe00;
			16'hb581: y = 16'hfe00;
			16'hb582: y = 16'hfe00;
			16'hb583: y = 16'hfe00;
			16'hb584: y = 16'hfe00;
			16'hb585: y = 16'hfe00;
			16'hb586: y = 16'hfe00;
			16'hb587: y = 16'hfe00;
			16'hb588: y = 16'hfe00;
			16'hb589: y = 16'hfe00;
			16'hb58a: y = 16'hfe00;
			16'hb58b: y = 16'hfe00;
			16'hb58c: y = 16'hfe00;
			16'hb58d: y = 16'hfe00;
			16'hb58e: y = 16'hfe00;
			16'hb58f: y = 16'hfe00;
			16'hb590: y = 16'hfe00;
			16'hb591: y = 16'hfe00;
			16'hb592: y = 16'hfe00;
			16'hb593: y = 16'hfe00;
			16'hb594: y = 16'hfe00;
			16'hb595: y = 16'hfe00;
			16'hb596: y = 16'hfe00;
			16'hb597: y = 16'hfe00;
			16'hb598: y = 16'hfe00;
			16'hb599: y = 16'hfe00;
			16'hb59a: y = 16'hfe00;
			16'hb59b: y = 16'hfe00;
			16'hb59c: y = 16'hfe00;
			16'hb59d: y = 16'hfe00;
			16'hb59e: y = 16'hfe00;
			16'hb59f: y = 16'hfe00;
			16'hb5a0: y = 16'hfe00;
			16'hb5a1: y = 16'hfe00;
			16'hb5a2: y = 16'hfe00;
			16'hb5a3: y = 16'hfe00;
			16'hb5a4: y = 16'hfe00;
			16'hb5a5: y = 16'hfe00;
			16'hb5a6: y = 16'hfe00;
			16'hb5a7: y = 16'hfe00;
			16'hb5a8: y = 16'hfe00;
			16'hb5a9: y = 16'hfe00;
			16'hb5aa: y = 16'hfe00;
			16'hb5ab: y = 16'hfe00;
			16'hb5ac: y = 16'hfe00;
			16'hb5ad: y = 16'hfe00;
			16'hb5ae: y = 16'hfe00;
			16'hb5af: y = 16'hfe00;
			16'hb5b0: y = 16'hfe00;
			16'hb5b1: y = 16'hfe00;
			16'hb5b2: y = 16'hfe00;
			16'hb5b3: y = 16'hfe00;
			16'hb5b4: y = 16'hfe00;
			16'hb5b5: y = 16'hfe00;
			16'hb5b6: y = 16'hfe00;
			16'hb5b7: y = 16'hfe00;
			16'hb5b8: y = 16'hfe00;
			16'hb5b9: y = 16'hfe00;
			16'hb5ba: y = 16'hfe00;
			16'hb5bb: y = 16'hfe00;
			16'hb5bc: y = 16'hfe00;
			16'hb5bd: y = 16'hfe00;
			16'hb5be: y = 16'hfe00;
			16'hb5bf: y = 16'hfe00;
			16'hb5c0: y = 16'hfe00;
			16'hb5c1: y = 16'hfe00;
			16'hb5c2: y = 16'hfe00;
			16'hb5c3: y = 16'hfe00;
			16'hb5c4: y = 16'hfe00;
			16'hb5c5: y = 16'hfe00;
			16'hb5c6: y = 16'hfe00;
			16'hb5c7: y = 16'hfe00;
			16'hb5c8: y = 16'hfe00;
			16'hb5c9: y = 16'hfe00;
			16'hb5ca: y = 16'hfe00;
			16'hb5cb: y = 16'hfe00;
			16'hb5cc: y = 16'hfe00;
			16'hb5cd: y = 16'hfe00;
			16'hb5ce: y = 16'hfe00;
			16'hb5cf: y = 16'hfe00;
			16'hb5d0: y = 16'hfe00;
			16'hb5d1: y = 16'hfe00;
			16'hb5d2: y = 16'hfe00;
			16'hb5d3: y = 16'hfe00;
			16'hb5d4: y = 16'hfe00;
			16'hb5d5: y = 16'hfe00;
			16'hb5d6: y = 16'hfe00;
			16'hb5d7: y = 16'hfe00;
			16'hb5d8: y = 16'hfe00;
			16'hb5d9: y = 16'hfe00;
			16'hb5da: y = 16'hfe00;
			16'hb5db: y = 16'hfe00;
			16'hb5dc: y = 16'hfe00;
			16'hb5dd: y = 16'hfe00;
			16'hb5de: y = 16'hfe00;
			16'hb5df: y = 16'hfe00;
			16'hb5e0: y = 16'hfe00;
			16'hb5e1: y = 16'hfe00;
			16'hb5e2: y = 16'hfe00;
			16'hb5e3: y = 16'hfe00;
			16'hb5e4: y = 16'hfe00;
			16'hb5e5: y = 16'hfe00;
			16'hb5e6: y = 16'hfe00;
			16'hb5e7: y = 16'hfe00;
			16'hb5e8: y = 16'hfe00;
			16'hb5e9: y = 16'hfe00;
			16'hb5ea: y = 16'hfe00;
			16'hb5eb: y = 16'hfe00;
			16'hb5ec: y = 16'hfe00;
			16'hb5ed: y = 16'hfe00;
			16'hb5ee: y = 16'hfe00;
			16'hb5ef: y = 16'hfe00;
			16'hb5f0: y = 16'hfe00;
			16'hb5f1: y = 16'hfe00;
			16'hb5f2: y = 16'hfe00;
			16'hb5f3: y = 16'hfe00;
			16'hb5f4: y = 16'hfe00;
			16'hb5f5: y = 16'hfe00;
			16'hb5f6: y = 16'hfe00;
			16'hb5f7: y = 16'hfe00;
			16'hb5f8: y = 16'hfe00;
			16'hb5f9: y = 16'hfe00;
			16'hb5fa: y = 16'hfe00;
			16'hb5fb: y = 16'hfe00;
			16'hb5fc: y = 16'hfe00;
			16'hb5fd: y = 16'hfe00;
			16'hb5fe: y = 16'hfe00;
			16'hb5ff: y = 16'hfe00;
			16'hb600: y = 16'hfe00;
			16'hb601: y = 16'hfe00;
			16'hb602: y = 16'hfe00;
			16'hb603: y = 16'hfe00;
			16'hb604: y = 16'hfe00;
			16'hb605: y = 16'hfe00;
			16'hb606: y = 16'hfe00;
			16'hb607: y = 16'hfe00;
			16'hb608: y = 16'hfe00;
			16'hb609: y = 16'hfe00;
			16'hb60a: y = 16'hfe00;
			16'hb60b: y = 16'hfe00;
			16'hb60c: y = 16'hfe00;
			16'hb60d: y = 16'hfe00;
			16'hb60e: y = 16'hfe00;
			16'hb60f: y = 16'hfe00;
			16'hb610: y = 16'hfe00;
			16'hb611: y = 16'hfe00;
			16'hb612: y = 16'hfe00;
			16'hb613: y = 16'hfe00;
			16'hb614: y = 16'hfe00;
			16'hb615: y = 16'hfe00;
			16'hb616: y = 16'hfe00;
			16'hb617: y = 16'hfe00;
			16'hb618: y = 16'hfe00;
			16'hb619: y = 16'hfe00;
			16'hb61a: y = 16'hfe00;
			16'hb61b: y = 16'hfe00;
			16'hb61c: y = 16'hfe00;
			16'hb61d: y = 16'hfe00;
			16'hb61e: y = 16'hfe00;
			16'hb61f: y = 16'hfe00;
			16'hb620: y = 16'hfe00;
			16'hb621: y = 16'hfe00;
			16'hb622: y = 16'hfe00;
			16'hb623: y = 16'hfe00;
			16'hb624: y = 16'hfe00;
			16'hb625: y = 16'hfe00;
			16'hb626: y = 16'hfe00;
			16'hb627: y = 16'hfe00;
			16'hb628: y = 16'hfe00;
			16'hb629: y = 16'hfe00;
			16'hb62a: y = 16'hfe00;
			16'hb62b: y = 16'hfe00;
			16'hb62c: y = 16'hfe00;
			16'hb62d: y = 16'hfe00;
			16'hb62e: y = 16'hfe00;
			16'hb62f: y = 16'hfe00;
			16'hb630: y = 16'hfe00;
			16'hb631: y = 16'hfe00;
			16'hb632: y = 16'hfe00;
			16'hb633: y = 16'hfe00;
			16'hb634: y = 16'hfe00;
			16'hb635: y = 16'hfe00;
			16'hb636: y = 16'hfe00;
			16'hb637: y = 16'hfe00;
			16'hb638: y = 16'hfe00;
			16'hb639: y = 16'hfe00;
			16'hb63a: y = 16'hfe00;
			16'hb63b: y = 16'hfe00;
			16'hb63c: y = 16'hfe00;
			16'hb63d: y = 16'hfe00;
			16'hb63e: y = 16'hfe00;
			16'hb63f: y = 16'hfe00;
			16'hb640: y = 16'hfe00;
			16'hb641: y = 16'hfe00;
			16'hb642: y = 16'hfe00;
			16'hb643: y = 16'hfe00;
			16'hb644: y = 16'hfe00;
			16'hb645: y = 16'hfe00;
			16'hb646: y = 16'hfe00;
			16'hb647: y = 16'hfe00;
			16'hb648: y = 16'hfe00;
			16'hb649: y = 16'hfe00;
			16'hb64a: y = 16'hfe00;
			16'hb64b: y = 16'hfe00;
			16'hb64c: y = 16'hfe00;
			16'hb64d: y = 16'hfe00;
			16'hb64e: y = 16'hfe00;
			16'hb64f: y = 16'hfe00;
			16'hb650: y = 16'hfe00;
			16'hb651: y = 16'hfe00;
			16'hb652: y = 16'hfe00;
			16'hb653: y = 16'hfe00;
			16'hb654: y = 16'hfe00;
			16'hb655: y = 16'hfe00;
			16'hb656: y = 16'hfe00;
			16'hb657: y = 16'hfe00;
			16'hb658: y = 16'hfe00;
			16'hb659: y = 16'hfe00;
			16'hb65a: y = 16'hfe00;
			16'hb65b: y = 16'hfe00;
			16'hb65c: y = 16'hfe00;
			16'hb65d: y = 16'hfe00;
			16'hb65e: y = 16'hfe00;
			16'hb65f: y = 16'hfe00;
			16'hb660: y = 16'hfe00;
			16'hb661: y = 16'hfe00;
			16'hb662: y = 16'hfe00;
			16'hb663: y = 16'hfe00;
			16'hb664: y = 16'hfe00;
			16'hb665: y = 16'hfe00;
			16'hb666: y = 16'hfe00;
			16'hb667: y = 16'hfe00;
			16'hb668: y = 16'hfe00;
			16'hb669: y = 16'hfe00;
			16'hb66a: y = 16'hfe00;
			16'hb66b: y = 16'hfe00;
			16'hb66c: y = 16'hfe00;
			16'hb66d: y = 16'hfe00;
			16'hb66e: y = 16'hfe00;
			16'hb66f: y = 16'hfe00;
			16'hb670: y = 16'hfe00;
			16'hb671: y = 16'hfe00;
			16'hb672: y = 16'hfe00;
			16'hb673: y = 16'hfe00;
			16'hb674: y = 16'hfe00;
			16'hb675: y = 16'hfe00;
			16'hb676: y = 16'hfe00;
			16'hb677: y = 16'hfe00;
			16'hb678: y = 16'hfe00;
			16'hb679: y = 16'hfe00;
			16'hb67a: y = 16'hfe00;
			16'hb67b: y = 16'hfe00;
			16'hb67c: y = 16'hfe00;
			16'hb67d: y = 16'hfe00;
			16'hb67e: y = 16'hfe00;
			16'hb67f: y = 16'hfe00;
			16'hb680: y = 16'hfe00;
			16'hb681: y = 16'hfe00;
			16'hb682: y = 16'hfe00;
			16'hb683: y = 16'hfe00;
			16'hb684: y = 16'hfe00;
			16'hb685: y = 16'hfe00;
			16'hb686: y = 16'hfe00;
			16'hb687: y = 16'hfe00;
			16'hb688: y = 16'hfe00;
			16'hb689: y = 16'hfe00;
			16'hb68a: y = 16'hfe00;
			16'hb68b: y = 16'hfe00;
			16'hb68c: y = 16'hfe00;
			16'hb68d: y = 16'hfe00;
			16'hb68e: y = 16'hfe00;
			16'hb68f: y = 16'hfe00;
			16'hb690: y = 16'hfe00;
			16'hb691: y = 16'hfe00;
			16'hb692: y = 16'hfe00;
			16'hb693: y = 16'hfe00;
			16'hb694: y = 16'hfe00;
			16'hb695: y = 16'hfe00;
			16'hb696: y = 16'hfe00;
			16'hb697: y = 16'hfe00;
			16'hb698: y = 16'hfe00;
			16'hb699: y = 16'hfe00;
			16'hb69a: y = 16'hfe00;
			16'hb69b: y = 16'hfe00;
			16'hb69c: y = 16'hfe00;
			16'hb69d: y = 16'hfe00;
			16'hb69e: y = 16'hfe00;
			16'hb69f: y = 16'hfe00;
			16'hb6a0: y = 16'hfe00;
			16'hb6a1: y = 16'hfe00;
			16'hb6a2: y = 16'hfe00;
			16'hb6a3: y = 16'hfe00;
			16'hb6a4: y = 16'hfe00;
			16'hb6a5: y = 16'hfe00;
			16'hb6a6: y = 16'hfe00;
			16'hb6a7: y = 16'hfe00;
			16'hb6a8: y = 16'hfe00;
			16'hb6a9: y = 16'hfe00;
			16'hb6aa: y = 16'hfe00;
			16'hb6ab: y = 16'hfe00;
			16'hb6ac: y = 16'hfe00;
			16'hb6ad: y = 16'hfe00;
			16'hb6ae: y = 16'hfe00;
			16'hb6af: y = 16'hfe00;
			16'hb6b0: y = 16'hfe00;
			16'hb6b1: y = 16'hfe00;
			16'hb6b2: y = 16'hfe00;
			16'hb6b3: y = 16'hfe00;
			16'hb6b4: y = 16'hfe00;
			16'hb6b5: y = 16'hfe00;
			16'hb6b6: y = 16'hfe00;
			16'hb6b7: y = 16'hfe00;
			16'hb6b8: y = 16'hfe00;
			16'hb6b9: y = 16'hfe00;
			16'hb6ba: y = 16'hfe00;
			16'hb6bb: y = 16'hfe00;
			16'hb6bc: y = 16'hfe00;
			16'hb6bd: y = 16'hfe00;
			16'hb6be: y = 16'hfe00;
			16'hb6bf: y = 16'hfe00;
			16'hb6c0: y = 16'hfe00;
			16'hb6c1: y = 16'hfe00;
			16'hb6c2: y = 16'hfe00;
			16'hb6c3: y = 16'hfe00;
			16'hb6c4: y = 16'hfe00;
			16'hb6c5: y = 16'hfe00;
			16'hb6c6: y = 16'hfe00;
			16'hb6c7: y = 16'hfe00;
			16'hb6c8: y = 16'hfe00;
			16'hb6c9: y = 16'hfe00;
			16'hb6ca: y = 16'hfe00;
			16'hb6cb: y = 16'hfe00;
			16'hb6cc: y = 16'hfe00;
			16'hb6cd: y = 16'hfe00;
			16'hb6ce: y = 16'hfe00;
			16'hb6cf: y = 16'hfe00;
			16'hb6d0: y = 16'hfe00;
			16'hb6d1: y = 16'hfe00;
			16'hb6d2: y = 16'hfe00;
			16'hb6d3: y = 16'hfe00;
			16'hb6d4: y = 16'hfe00;
			16'hb6d5: y = 16'hfe00;
			16'hb6d6: y = 16'hfe00;
			16'hb6d7: y = 16'hfe00;
			16'hb6d8: y = 16'hfe00;
			16'hb6d9: y = 16'hfe00;
			16'hb6da: y = 16'hfe00;
			16'hb6db: y = 16'hfe00;
			16'hb6dc: y = 16'hfe00;
			16'hb6dd: y = 16'hfe00;
			16'hb6de: y = 16'hfe00;
			16'hb6df: y = 16'hfe00;
			16'hb6e0: y = 16'hfe00;
			16'hb6e1: y = 16'hfe00;
			16'hb6e2: y = 16'hfe00;
			16'hb6e3: y = 16'hfe00;
			16'hb6e4: y = 16'hfe00;
			16'hb6e5: y = 16'hfe00;
			16'hb6e6: y = 16'hfe00;
			16'hb6e7: y = 16'hfe00;
			16'hb6e8: y = 16'hfe00;
			16'hb6e9: y = 16'hfe00;
			16'hb6ea: y = 16'hfe00;
			16'hb6eb: y = 16'hfe00;
			16'hb6ec: y = 16'hfe00;
			16'hb6ed: y = 16'hfe00;
			16'hb6ee: y = 16'hfe00;
			16'hb6ef: y = 16'hfe00;
			16'hb6f0: y = 16'hfe00;
			16'hb6f1: y = 16'hfe00;
			16'hb6f2: y = 16'hfe00;
			16'hb6f3: y = 16'hfe00;
			16'hb6f4: y = 16'hfe00;
			16'hb6f5: y = 16'hfe00;
			16'hb6f6: y = 16'hfe00;
			16'hb6f7: y = 16'hfe00;
			16'hb6f8: y = 16'hfe00;
			16'hb6f9: y = 16'hfe00;
			16'hb6fa: y = 16'hfe00;
			16'hb6fb: y = 16'hfe00;
			16'hb6fc: y = 16'hfe00;
			16'hb6fd: y = 16'hfe00;
			16'hb6fe: y = 16'hfe00;
			16'hb6ff: y = 16'hfe00;
			16'hb700: y = 16'hfe00;
			16'hb701: y = 16'hfe00;
			16'hb702: y = 16'hfe00;
			16'hb703: y = 16'hfe00;
			16'hb704: y = 16'hfe00;
			16'hb705: y = 16'hfe00;
			16'hb706: y = 16'hfe00;
			16'hb707: y = 16'hfe00;
			16'hb708: y = 16'hfe00;
			16'hb709: y = 16'hfe00;
			16'hb70a: y = 16'hfe00;
			16'hb70b: y = 16'hfe00;
			16'hb70c: y = 16'hfe00;
			16'hb70d: y = 16'hfe00;
			16'hb70e: y = 16'hfe00;
			16'hb70f: y = 16'hfe00;
			16'hb710: y = 16'hfe00;
			16'hb711: y = 16'hfe00;
			16'hb712: y = 16'hfe00;
			16'hb713: y = 16'hfe00;
			16'hb714: y = 16'hfe00;
			16'hb715: y = 16'hfe00;
			16'hb716: y = 16'hfe00;
			16'hb717: y = 16'hfe00;
			16'hb718: y = 16'hfe00;
			16'hb719: y = 16'hfe00;
			16'hb71a: y = 16'hfe00;
			16'hb71b: y = 16'hfe00;
			16'hb71c: y = 16'hfe00;
			16'hb71d: y = 16'hfe00;
			16'hb71e: y = 16'hfe00;
			16'hb71f: y = 16'hfe00;
			16'hb720: y = 16'hfe00;
			16'hb721: y = 16'hfe00;
			16'hb722: y = 16'hfe00;
			16'hb723: y = 16'hfe00;
			16'hb724: y = 16'hfe00;
			16'hb725: y = 16'hfe00;
			16'hb726: y = 16'hfe00;
			16'hb727: y = 16'hfe00;
			16'hb728: y = 16'hfe00;
			16'hb729: y = 16'hfe00;
			16'hb72a: y = 16'hfe00;
			16'hb72b: y = 16'hfe00;
			16'hb72c: y = 16'hfe00;
			16'hb72d: y = 16'hfe00;
			16'hb72e: y = 16'hfe00;
			16'hb72f: y = 16'hfe00;
			16'hb730: y = 16'hfe00;
			16'hb731: y = 16'hfe00;
			16'hb732: y = 16'hfe00;
			16'hb733: y = 16'hfe00;
			16'hb734: y = 16'hfe00;
			16'hb735: y = 16'hfe00;
			16'hb736: y = 16'hfe00;
			16'hb737: y = 16'hfe00;
			16'hb738: y = 16'hfe00;
			16'hb739: y = 16'hfe00;
			16'hb73a: y = 16'hfe00;
			16'hb73b: y = 16'hfe00;
			16'hb73c: y = 16'hfe00;
			16'hb73d: y = 16'hfe00;
			16'hb73e: y = 16'hfe00;
			16'hb73f: y = 16'hfe00;
			16'hb740: y = 16'hfe00;
			16'hb741: y = 16'hfe00;
			16'hb742: y = 16'hfe00;
			16'hb743: y = 16'hfe00;
			16'hb744: y = 16'hfe00;
			16'hb745: y = 16'hfe00;
			16'hb746: y = 16'hfe00;
			16'hb747: y = 16'hfe00;
			16'hb748: y = 16'hfe00;
			16'hb749: y = 16'hfe00;
			16'hb74a: y = 16'hfe00;
			16'hb74b: y = 16'hfe00;
			16'hb74c: y = 16'hfe00;
			16'hb74d: y = 16'hfe00;
			16'hb74e: y = 16'hfe00;
			16'hb74f: y = 16'hfe00;
			16'hb750: y = 16'hfe00;
			16'hb751: y = 16'hfe00;
			16'hb752: y = 16'hfe00;
			16'hb753: y = 16'hfe00;
			16'hb754: y = 16'hfe00;
			16'hb755: y = 16'hfe00;
			16'hb756: y = 16'hfe00;
			16'hb757: y = 16'hfe00;
			16'hb758: y = 16'hfe00;
			16'hb759: y = 16'hfe00;
			16'hb75a: y = 16'hfe00;
			16'hb75b: y = 16'hfe00;
			16'hb75c: y = 16'hfe00;
			16'hb75d: y = 16'hfe00;
			16'hb75e: y = 16'hfe00;
			16'hb75f: y = 16'hfe00;
			16'hb760: y = 16'hfe00;
			16'hb761: y = 16'hfe00;
			16'hb762: y = 16'hfe00;
			16'hb763: y = 16'hfe00;
			16'hb764: y = 16'hfe00;
			16'hb765: y = 16'hfe00;
			16'hb766: y = 16'hfe00;
			16'hb767: y = 16'hfe00;
			16'hb768: y = 16'hfe00;
			16'hb769: y = 16'hfe00;
			16'hb76a: y = 16'hfe00;
			16'hb76b: y = 16'hfe00;
			16'hb76c: y = 16'hfe00;
			16'hb76d: y = 16'hfe00;
			16'hb76e: y = 16'hfe00;
			16'hb76f: y = 16'hfe00;
			16'hb770: y = 16'hfe00;
			16'hb771: y = 16'hfe00;
			16'hb772: y = 16'hfe00;
			16'hb773: y = 16'hfe00;
			16'hb774: y = 16'hfe00;
			16'hb775: y = 16'hfe00;
			16'hb776: y = 16'hfe00;
			16'hb777: y = 16'hfe00;
			16'hb778: y = 16'hfe00;
			16'hb779: y = 16'hfe00;
			16'hb77a: y = 16'hfe00;
			16'hb77b: y = 16'hfe00;
			16'hb77c: y = 16'hfe00;
			16'hb77d: y = 16'hfe00;
			16'hb77e: y = 16'hfe00;
			16'hb77f: y = 16'hfe00;
			16'hb780: y = 16'hfe00;
			16'hb781: y = 16'hfe00;
			16'hb782: y = 16'hfe00;
			16'hb783: y = 16'hfe00;
			16'hb784: y = 16'hfe00;
			16'hb785: y = 16'hfe00;
			16'hb786: y = 16'hfe00;
			16'hb787: y = 16'hfe00;
			16'hb788: y = 16'hfe00;
			16'hb789: y = 16'hfe00;
			16'hb78a: y = 16'hfe00;
			16'hb78b: y = 16'hfe00;
			16'hb78c: y = 16'hfe00;
			16'hb78d: y = 16'hfe00;
			16'hb78e: y = 16'hfe00;
			16'hb78f: y = 16'hfe00;
			16'hb790: y = 16'hfe00;
			16'hb791: y = 16'hfe00;
			16'hb792: y = 16'hfe00;
			16'hb793: y = 16'hfe00;
			16'hb794: y = 16'hfe00;
			16'hb795: y = 16'hfe00;
			16'hb796: y = 16'hfe00;
			16'hb797: y = 16'hfe00;
			16'hb798: y = 16'hfe00;
			16'hb799: y = 16'hfe00;
			16'hb79a: y = 16'hfe00;
			16'hb79b: y = 16'hfe00;
			16'hb79c: y = 16'hfe00;
			16'hb79d: y = 16'hfe00;
			16'hb79e: y = 16'hfe00;
			16'hb79f: y = 16'hfe00;
			16'hb7a0: y = 16'hfe00;
			16'hb7a1: y = 16'hfe00;
			16'hb7a2: y = 16'hfe00;
			16'hb7a3: y = 16'hfe00;
			16'hb7a4: y = 16'hfe00;
			16'hb7a5: y = 16'hfe00;
			16'hb7a6: y = 16'hfe00;
			16'hb7a7: y = 16'hfe00;
			16'hb7a8: y = 16'hfe00;
			16'hb7a9: y = 16'hfe00;
			16'hb7aa: y = 16'hfe00;
			16'hb7ab: y = 16'hfe00;
			16'hb7ac: y = 16'hfe00;
			16'hb7ad: y = 16'hfe00;
			16'hb7ae: y = 16'hfe00;
			16'hb7af: y = 16'hfe00;
			16'hb7b0: y = 16'hfe00;
			16'hb7b1: y = 16'hfe00;
			16'hb7b2: y = 16'hfe00;
			16'hb7b3: y = 16'hfe00;
			16'hb7b4: y = 16'hfe00;
			16'hb7b5: y = 16'hfe00;
			16'hb7b6: y = 16'hfe00;
			16'hb7b7: y = 16'hfe00;
			16'hb7b8: y = 16'hfe00;
			16'hb7b9: y = 16'hfe00;
			16'hb7ba: y = 16'hfe00;
			16'hb7bb: y = 16'hfe00;
			16'hb7bc: y = 16'hfe00;
			16'hb7bd: y = 16'hfe00;
			16'hb7be: y = 16'hfe00;
			16'hb7bf: y = 16'hfe00;
			16'hb7c0: y = 16'hfe00;
			16'hb7c1: y = 16'hfe00;
			16'hb7c2: y = 16'hfe00;
			16'hb7c3: y = 16'hfe00;
			16'hb7c4: y = 16'hfe00;
			16'hb7c5: y = 16'hfe00;
			16'hb7c6: y = 16'hfe00;
			16'hb7c7: y = 16'hfe00;
			16'hb7c8: y = 16'hfe00;
			16'hb7c9: y = 16'hfe00;
			16'hb7ca: y = 16'hfe00;
			16'hb7cb: y = 16'hfe00;
			16'hb7cc: y = 16'hfe00;
			16'hb7cd: y = 16'hfe00;
			16'hb7ce: y = 16'hfe00;
			16'hb7cf: y = 16'hfe00;
			16'hb7d0: y = 16'hfe00;
			16'hb7d1: y = 16'hfe00;
			16'hb7d2: y = 16'hfe00;
			16'hb7d3: y = 16'hfe00;
			16'hb7d4: y = 16'hfe00;
			16'hb7d5: y = 16'hfe00;
			16'hb7d6: y = 16'hfe00;
			16'hb7d7: y = 16'hfe00;
			16'hb7d8: y = 16'hfe00;
			16'hb7d9: y = 16'hfe00;
			16'hb7da: y = 16'hfe00;
			16'hb7db: y = 16'hfe00;
			16'hb7dc: y = 16'hfe00;
			16'hb7dd: y = 16'hfe00;
			16'hb7de: y = 16'hfe00;
			16'hb7df: y = 16'hfe00;
			16'hb7e0: y = 16'hfe00;
			16'hb7e1: y = 16'hfe00;
			16'hb7e2: y = 16'hfe00;
			16'hb7e3: y = 16'hfe00;
			16'hb7e4: y = 16'hfe00;
			16'hb7e5: y = 16'hfe00;
			16'hb7e6: y = 16'hfe00;
			16'hb7e7: y = 16'hfe00;
			16'hb7e8: y = 16'hfe00;
			16'hb7e9: y = 16'hfe00;
			16'hb7ea: y = 16'hfe00;
			16'hb7eb: y = 16'hfe00;
			16'hb7ec: y = 16'hfe00;
			16'hb7ed: y = 16'hfe00;
			16'hb7ee: y = 16'hfe00;
			16'hb7ef: y = 16'hfe00;
			16'hb7f0: y = 16'hfe00;
			16'hb7f1: y = 16'hfe00;
			16'hb7f2: y = 16'hfe00;
			16'hb7f3: y = 16'hfe00;
			16'hb7f4: y = 16'hfe00;
			16'hb7f5: y = 16'hfe00;
			16'hb7f6: y = 16'hfe00;
			16'hb7f7: y = 16'hfe00;
			16'hb7f8: y = 16'hfe00;
			16'hb7f9: y = 16'hfe00;
			16'hb7fa: y = 16'hfe00;
			16'hb7fb: y = 16'hfe00;
			16'hb7fc: y = 16'hfe00;
			16'hb7fd: y = 16'hfe00;
			16'hb7fe: y = 16'hfe00;
			16'hb7ff: y = 16'hfe00;
			16'hb800: y = 16'hfe00;
			16'hb801: y = 16'hfe00;
			16'hb802: y = 16'hfe00;
			16'hb803: y = 16'hfe00;
			16'hb804: y = 16'hfe00;
			16'hb805: y = 16'hfe00;
			16'hb806: y = 16'hfe00;
			16'hb807: y = 16'hfe00;
			16'hb808: y = 16'hfe00;
			16'hb809: y = 16'hfe00;
			16'hb80a: y = 16'hfe00;
			16'hb80b: y = 16'hfe00;
			16'hb80c: y = 16'hfe00;
			16'hb80d: y = 16'hfe00;
			16'hb80e: y = 16'hfe00;
			16'hb80f: y = 16'hfe00;
			16'hb810: y = 16'hfe00;
			16'hb811: y = 16'hfe00;
			16'hb812: y = 16'hfe00;
			16'hb813: y = 16'hfe00;
			16'hb814: y = 16'hfe00;
			16'hb815: y = 16'hfe00;
			16'hb816: y = 16'hfe00;
			16'hb817: y = 16'hfe00;
			16'hb818: y = 16'hfe00;
			16'hb819: y = 16'hfe00;
			16'hb81a: y = 16'hfe00;
			16'hb81b: y = 16'hfe00;
			16'hb81c: y = 16'hfe00;
			16'hb81d: y = 16'hfe00;
			16'hb81e: y = 16'hfe00;
			16'hb81f: y = 16'hfe00;
			16'hb820: y = 16'hfe00;
			16'hb821: y = 16'hfe00;
			16'hb822: y = 16'hfe00;
			16'hb823: y = 16'hfe00;
			16'hb824: y = 16'hfe00;
			16'hb825: y = 16'hfe00;
			16'hb826: y = 16'hfe00;
			16'hb827: y = 16'hfe00;
			16'hb828: y = 16'hfe00;
			16'hb829: y = 16'hfe00;
			16'hb82a: y = 16'hfe00;
			16'hb82b: y = 16'hfe00;
			16'hb82c: y = 16'hfe00;
			16'hb82d: y = 16'hfe00;
			16'hb82e: y = 16'hfe00;
			16'hb82f: y = 16'hfe00;
			16'hb830: y = 16'hfe00;
			16'hb831: y = 16'hfe00;
			16'hb832: y = 16'hfe00;
			16'hb833: y = 16'hfe00;
			16'hb834: y = 16'hfe00;
			16'hb835: y = 16'hfe00;
			16'hb836: y = 16'hfe00;
			16'hb837: y = 16'hfe00;
			16'hb838: y = 16'hfe00;
			16'hb839: y = 16'hfe00;
			16'hb83a: y = 16'hfe00;
			16'hb83b: y = 16'hfe00;
			16'hb83c: y = 16'hfe00;
			16'hb83d: y = 16'hfe00;
			16'hb83e: y = 16'hfe00;
			16'hb83f: y = 16'hfe00;
			16'hb840: y = 16'hfe00;
			16'hb841: y = 16'hfe00;
			16'hb842: y = 16'hfe00;
			16'hb843: y = 16'hfe00;
			16'hb844: y = 16'hfe00;
			16'hb845: y = 16'hfe00;
			16'hb846: y = 16'hfe00;
			16'hb847: y = 16'hfe00;
			16'hb848: y = 16'hfe00;
			16'hb849: y = 16'hfe00;
			16'hb84a: y = 16'hfe00;
			16'hb84b: y = 16'hfe00;
			16'hb84c: y = 16'hfe00;
			16'hb84d: y = 16'hfe00;
			16'hb84e: y = 16'hfe00;
			16'hb84f: y = 16'hfe00;
			16'hb850: y = 16'hfe00;
			16'hb851: y = 16'hfe00;
			16'hb852: y = 16'hfe00;
			16'hb853: y = 16'hfe00;
			16'hb854: y = 16'hfe00;
			16'hb855: y = 16'hfe00;
			16'hb856: y = 16'hfe00;
			16'hb857: y = 16'hfe00;
			16'hb858: y = 16'hfe00;
			16'hb859: y = 16'hfe00;
			16'hb85a: y = 16'hfe00;
			16'hb85b: y = 16'hfe00;
			16'hb85c: y = 16'hfe00;
			16'hb85d: y = 16'hfe00;
			16'hb85e: y = 16'hfe00;
			16'hb85f: y = 16'hfe00;
			16'hb860: y = 16'hfe00;
			16'hb861: y = 16'hfe00;
			16'hb862: y = 16'hfe00;
			16'hb863: y = 16'hfe00;
			16'hb864: y = 16'hfe00;
			16'hb865: y = 16'hfe00;
			16'hb866: y = 16'hfe00;
			16'hb867: y = 16'hfe00;
			16'hb868: y = 16'hfe00;
			16'hb869: y = 16'hfe00;
			16'hb86a: y = 16'hfe00;
			16'hb86b: y = 16'hfe00;
			16'hb86c: y = 16'hfe00;
			16'hb86d: y = 16'hfe00;
			16'hb86e: y = 16'hfe00;
			16'hb86f: y = 16'hfe00;
			16'hb870: y = 16'hfe00;
			16'hb871: y = 16'hfe00;
			16'hb872: y = 16'hfe00;
			16'hb873: y = 16'hfe00;
			16'hb874: y = 16'hfe00;
			16'hb875: y = 16'hfe00;
			16'hb876: y = 16'hfe00;
			16'hb877: y = 16'hfe00;
			16'hb878: y = 16'hfe00;
			16'hb879: y = 16'hfe00;
			16'hb87a: y = 16'hfe00;
			16'hb87b: y = 16'hfe00;
			16'hb87c: y = 16'hfe00;
			16'hb87d: y = 16'hfe00;
			16'hb87e: y = 16'hfe00;
			16'hb87f: y = 16'hfe00;
			16'hb880: y = 16'hfe00;
			16'hb881: y = 16'hfe00;
			16'hb882: y = 16'hfe00;
			16'hb883: y = 16'hfe00;
			16'hb884: y = 16'hfe00;
			16'hb885: y = 16'hfe00;
			16'hb886: y = 16'hfe00;
			16'hb887: y = 16'hfe00;
			16'hb888: y = 16'hfe00;
			16'hb889: y = 16'hfe00;
			16'hb88a: y = 16'hfe00;
			16'hb88b: y = 16'hfe00;
			16'hb88c: y = 16'hfe00;
			16'hb88d: y = 16'hfe00;
			16'hb88e: y = 16'hfe00;
			16'hb88f: y = 16'hfe00;
			16'hb890: y = 16'hfe00;
			16'hb891: y = 16'hfe00;
			16'hb892: y = 16'hfe00;
			16'hb893: y = 16'hfe00;
			16'hb894: y = 16'hfe00;
			16'hb895: y = 16'hfe00;
			16'hb896: y = 16'hfe00;
			16'hb897: y = 16'hfe00;
			16'hb898: y = 16'hfe00;
			16'hb899: y = 16'hfe00;
			16'hb89a: y = 16'hfe00;
			16'hb89b: y = 16'hfe00;
			16'hb89c: y = 16'hfe00;
			16'hb89d: y = 16'hfe00;
			16'hb89e: y = 16'hfe00;
			16'hb89f: y = 16'hfe00;
			16'hb8a0: y = 16'hfe00;
			16'hb8a1: y = 16'hfe00;
			16'hb8a2: y = 16'hfe00;
			16'hb8a3: y = 16'hfe00;
			16'hb8a4: y = 16'hfe00;
			16'hb8a5: y = 16'hfe00;
			16'hb8a6: y = 16'hfe00;
			16'hb8a7: y = 16'hfe00;
			16'hb8a8: y = 16'hfe00;
			16'hb8a9: y = 16'hfe00;
			16'hb8aa: y = 16'hfe00;
			16'hb8ab: y = 16'hfe00;
			16'hb8ac: y = 16'hfe00;
			16'hb8ad: y = 16'hfe00;
			16'hb8ae: y = 16'hfe00;
			16'hb8af: y = 16'hfe00;
			16'hb8b0: y = 16'hfe00;
			16'hb8b1: y = 16'hfe00;
			16'hb8b2: y = 16'hfe00;
			16'hb8b3: y = 16'hfe00;
			16'hb8b4: y = 16'hfe00;
			16'hb8b5: y = 16'hfe00;
			16'hb8b6: y = 16'hfe00;
			16'hb8b7: y = 16'hfe00;
			16'hb8b8: y = 16'hfe00;
			16'hb8b9: y = 16'hfe00;
			16'hb8ba: y = 16'hfe00;
			16'hb8bb: y = 16'hfe00;
			16'hb8bc: y = 16'hfe00;
			16'hb8bd: y = 16'hfe00;
			16'hb8be: y = 16'hfe00;
			16'hb8bf: y = 16'hfe00;
			16'hb8c0: y = 16'hfe00;
			16'hb8c1: y = 16'hfe00;
			16'hb8c2: y = 16'hfe00;
			16'hb8c3: y = 16'hfe00;
			16'hb8c4: y = 16'hfe00;
			16'hb8c5: y = 16'hfe00;
			16'hb8c6: y = 16'hfe00;
			16'hb8c7: y = 16'hfe00;
			16'hb8c8: y = 16'hfe00;
			16'hb8c9: y = 16'hfe00;
			16'hb8ca: y = 16'hfe00;
			16'hb8cb: y = 16'hfe00;
			16'hb8cc: y = 16'hfe00;
			16'hb8cd: y = 16'hfe00;
			16'hb8ce: y = 16'hfe00;
			16'hb8cf: y = 16'hfe00;
			16'hb8d0: y = 16'hfe00;
			16'hb8d1: y = 16'hfe00;
			16'hb8d2: y = 16'hfe00;
			16'hb8d3: y = 16'hfe00;
			16'hb8d4: y = 16'hfe00;
			16'hb8d5: y = 16'hfe00;
			16'hb8d6: y = 16'hfe00;
			16'hb8d7: y = 16'hfe00;
			16'hb8d8: y = 16'hfe00;
			16'hb8d9: y = 16'hfe00;
			16'hb8da: y = 16'hfe00;
			16'hb8db: y = 16'hfe00;
			16'hb8dc: y = 16'hfe00;
			16'hb8dd: y = 16'hfe00;
			16'hb8de: y = 16'hfe00;
			16'hb8df: y = 16'hfe00;
			16'hb8e0: y = 16'hfe00;
			16'hb8e1: y = 16'hfe00;
			16'hb8e2: y = 16'hfe00;
			16'hb8e3: y = 16'hfe00;
			16'hb8e4: y = 16'hfe00;
			16'hb8e5: y = 16'hfe00;
			16'hb8e6: y = 16'hfe00;
			16'hb8e7: y = 16'hfe00;
			16'hb8e8: y = 16'hfe00;
			16'hb8e9: y = 16'hfe00;
			16'hb8ea: y = 16'hfe00;
			16'hb8eb: y = 16'hfe00;
			16'hb8ec: y = 16'hfe00;
			16'hb8ed: y = 16'hfe00;
			16'hb8ee: y = 16'hfe00;
			16'hb8ef: y = 16'hfe00;
			16'hb8f0: y = 16'hfe00;
			16'hb8f1: y = 16'hfe00;
			16'hb8f2: y = 16'hfe00;
			16'hb8f3: y = 16'hfe00;
			16'hb8f4: y = 16'hfe00;
			16'hb8f5: y = 16'hfe00;
			16'hb8f6: y = 16'hfe00;
			16'hb8f7: y = 16'hfe00;
			16'hb8f8: y = 16'hfe00;
			16'hb8f9: y = 16'hfe00;
			16'hb8fa: y = 16'hfe00;
			16'hb8fb: y = 16'hfe00;
			16'hb8fc: y = 16'hfe00;
			16'hb8fd: y = 16'hfe00;
			16'hb8fe: y = 16'hfe00;
			16'hb8ff: y = 16'hfe00;
			16'hb900: y = 16'hfe00;
			16'hb901: y = 16'hfe00;
			16'hb902: y = 16'hfe00;
			16'hb903: y = 16'hfe00;
			16'hb904: y = 16'hfe00;
			16'hb905: y = 16'hfe00;
			16'hb906: y = 16'hfe00;
			16'hb907: y = 16'hfe00;
			16'hb908: y = 16'hfe00;
			16'hb909: y = 16'hfe00;
			16'hb90a: y = 16'hfe00;
			16'hb90b: y = 16'hfe00;
			16'hb90c: y = 16'hfe00;
			16'hb90d: y = 16'hfe00;
			16'hb90e: y = 16'hfe00;
			16'hb90f: y = 16'hfe00;
			16'hb910: y = 16'hfe00;
			16'hb911: y = 16'hfe00;
			16'hb912: y = 16'hfe00;
			16'hb913: y = 16'hfe00;
			16'hb914: y = 16'hfe00;
			16'hb915: y = 16'hfe00;
			16'hb916: y = 16'hfe00;
			16'hb917: y = 16'hfe00;
			16'hb918: y = 16'hfe00;
			16'hb919: y = 16'hfe00;
			16'hb91a: y = 16'hfe00;
			16'hb91b: y = 16'hfe00;
			16'hb91c: y = 16'hfe00;
			16'hb91d: y = 16'hfe00;
			16'hb91e: y = 16'hfe00;
			16'hb91f: y = 16'hfe00;
			16'hb920: y = 16'hfe00;
			16'hb921: y = 16'hfe00;
			16'hb922: y = 16'hfe00;
			16'hb923: y = 16'hfe00;
			16'hb924: y = 16'hfe00;
			16'hb925: y = 16'hfe00;
			16'hb926: y = 16'hfe00;
			16'hb927: y = 16'hfe00;
			16'hb928: y = 16'hfe00;
			16'hb929: y = 16'hfe00;
			16'hb92a: y = 16'hfe00;
			16'hb92b: y = 16'hfe00;
			16'hb92c: y = 16'hfe00;
			16'hb92d: y = 16'hfe00;
			16'hb92e: y = 16'hfe00;
			16'hb92f: y = 16'hfe00;
			16'hb930: y = 16'hfe00;
			16'hb931: y = 16'hfe00;
			16'hb932: y = 16'hfe00;
			16'hb933: y = 16'hfe00;
			16'hb934: y = 16'hfe00;
			16'hb935: y = 16'hfe00;
			16'hb936: y = 16'hfe00;
			16'hb937: y = 16'hfe00;
			16'hb938: y = 16'hfe00;
			16'hb939: y = 16'hfe00;
			16'hb93a: y = 16'hfe00;
			16'hb93b: y = 16'hfe00;
			16'hb93c: y = 16'hfe00;
			16'hb93d: y = 16'hfe00;
			16'hb93e: y = 16'hfe00;
			16'hb93f: y = 16'hfe00;
			16'hb940: y = 16'hfe00;
			16'hb941: y = 16'hfe00;
			16'hb942: y = 16'hfe00;
			16'hb943: y = 16'hfe00;
			16'hb944: y = 16'hfe00;
			16'hb945: y = 16'hfe00;
			16'hb946: y = 16'hfe00;
			16'hb947: y = 16'hfe00;
			16'hb948: y = 16'hfe00;
			16'hb949: y = 16'hfe00;
			16'hb94a: y = 16'hfe00;
			16'hb94b: y = 16'hfe00;
			16'hb94c: y = 16'hfe00;
			16'hb94d: y = 16'hfe00;
			16'hb94e: y = 16'hfe00;
			16'hb94f: y = 16'hfe00;
			16'hb950: y = 16'hfe00;
			16'hb951: y = 16'hfe00;
			16'hb952: y = 16'hfe00;
			16'hb953: y = 16'hfe00;
			16'hb954: y = 16'hfe00;
			16'hb955: y = 16'hfe00;
			16'hb956: y = 16'hfe00;
			16'hb957: y = 16'hfe00;
			16'hb958: y = 16'hfe00;
			16'hb959: y = 16'hfe00;
			16'hb95a: y = 16'hfe00;
			16'hb95b: y = 16'hfe00;
			16'hb95c: y = 16'hfe00;
			16'hb95d: y = 16'hfe00;
			16'hb95e: y = 16'hfe00;
			16'hb95f: y = 16'hfe00;
			16'hb960: y = 16'hfe00;
			16'hb961: y = 16'hfe00;
			16'hb962: y = 16'hfe00;
			16'hb963: y = 16'hfe00;
			16'hb964: y = 16'hfe00;
			16'hb965: y = 16'hfe00;
			16'hb966: y = 16'hfe00;
			16'hb967: y = 16'hfe00;
			16'hb968: y = 16'hfe00;
			16'hb969: y = 16'hfe00;
			16'hb96a: y = 16'hfe00;
			16'hb96b: y = 16'hfe00;
			16'hb96c: y = 16'hfe00;
			16'hb96d: y = 16'hfe00;
			16'hb96e: y = 16'hfe00;
			16'hb96f: y = 16'hfe00;
			16'hb970: y = 16'hfe00;
			16'hb971: y = 16'hfe00;
			16'hb972: y = 16'hfe00;
			16'hb973: y = 16'hfe00;
			16'hb974: y = 16'hfe00;
			16'hb975: y = 16'hfe00;
			16'hb976: y = 16'hfe00;
			16'hb977: y = 16'hfe00;
			16'hb978: y = 16'hfe00;
			16'hb979: y = 16'hfe00;
			16'hb97a: y = 16'hfe00;
			16'hb97b: y = 16'hfe00;
			16'hb97c: y = 16'hfe00;
			16'hb97d: y = 16'hfe00;
			16'hb97e: y = 16'hfe00;
			16'hb97f: y = 16'hfe00;
			16'hb980: y = 16'hfe00;
			16'hb981: y = 16'hfe00;
			16'hb982: y = 16'hfe00;
			16'hb983: y = 16'hfe00;
			16'hb984: y = 16'hfe00;
			16'hb985: y = 16'hfe00;
			16'hb986: y = 16'hfe00;
			16'hb987: y = 16'hfe00;
			16'hb988: y = 16'hfe00;
			16'hb989: y = 16'hfe00;
			16'hb98a: y = 16'hfe00;
			16'hb98b: y = 16'hfe00;
			16'hb98c: y = 16'hfe00;
			16'hb98d: y = 16'hfe00;
			16'hb98e: y = 16'hfe00;
			16'hb98f: y = 16'hfe00;
			16'hb990: y = 16'hfe00;
			16'hb991: y = 16'hfe00;
			16'hb992: y = 16'hfe00;
			16'hb993: y = 16'hfe00;
			16'hb994: y = 16'hfe00;
			16'hb995: y = 16'hfe00;
			16'hb996: y = 16'hfe00;
			16'hb997: y = 16'hfe00;
			16'hb998: y = 16'hfe00;
			16'hb999: y = 16'hfe00;
			16'hb99a: y = 16'hfe00;
			16'hb99b: y = 16'hfe00;
			16'hb99c: y = 16'hfe00;
			16'hb99d: y = 16'hfe00;
			16'hb99e: y = 16'hfe00;
			16'hb99f: y = 16'hfe00;
			16'hb9a0: y = 16'hfe00;
			16'hb9a1: y = 16'hfe00;
			16'hb9a2: y = 16'hfe00;
			16'hb9a3: y = 16'hfe00;
			16'hb9a4: y = 16'hfe00;
			16'hb9a5: y = 16'hfe00;
			16'hb9a6: y = 16'hfe00;
			16'hb9a7: y = 16'hfe00;
			16'hb9a8: y = 16'hfe00;
			16'hb9a9: y = 16'hfe00;
			16'hb9aa: y = 16'hfe00;
			16'hb9ab: y = 16'hfe00;
			16'hb9ac: y = 16'hfe00;
			16'hb9ad: y = 16'hfe00;
			16'hb9ae: y = 16'hfe00;
			16'hb9af: y = 16'hfe00;
			16'hb9b0: y = 16'hfe00;
			16'hb9b1: y = 16'hfe00;
			16'hb9b2: y = 16'hfe00;
			16'hb9b3: y = 16'hfe00;
			16'hb9b4: y = 16'hfe00;
			16'hb9b5: y = 16'hfe00;
			16'hb9b6: y = 16'hfe00;
			16'hb9b7: y = 16'hfe00;
			16'hb9b8: y = 16'hfe00;
			16'hb9b9: y = 16'hfe00;
			16'hb9ba: y = 16'hfe00;
			16'hb9bb: y = 16'hfe00;
			16'hb9bc: y = 16'hfe00;
			16'hb9bd: y = 16'hfe00;
			16'hb9be: y = 16'hfe00;
			16'hb9bf: y = 16'hfe00;
			16'hb9c0: y = 16'hfe00;
			16'hb9c1: y = 16'hfe00;
			16'hb9c2: y = 16'hfe00;
			16'hb9c3: y = 16'hfe00;
			16'hb9c4: y = 16'hfe00;
			16'hb9c5: y = 16'hfe00;
			16'hb9c6: y = 16'hfe00;
			16'hb9c7: y = 16'hfe00;
			16'hb9c8: y = 16'hfe00;
			16'hb9c9: y = 16'hfe00;
			16'hb9ca: y = 16'hfe00;
			16'hb9cb: y = 16'hfe00;
			16'hb9cc: y = 16'hfe00;
			16'hb9cd: y = 16'hfe00;
			16'hb9ce: y = 16'hfe00;
			16'hb9cf: y = 16'hfe00;
			16'hb9d0: y = 16'hfe00;
			16'hb9d1: y = 16'hfe00;
			16'hb9d2: y = 16'hfe00;
			16'hb9d3: y = 16'hfe00;
			16'hb9d4: y = 16'hfe00;
			16'hb9d5: y = 16'hfe00;
			16'hb9d6: y = 16'hfe00;
			16'hb9d7: y = 16'hfe00;
			16'hb9d8: y = 16'hfe00;
			16'hb9d9: y = 16'hfe00;
			16'hb9da: y = 16'hfe00;
			16'hb9db: y = 16'hfe00;
			16'hb9dc: y = 16'hfe00;
			16'hb9dd: y = 16'hfe00;
			16'hb9de: y = 16'hfe00;
			16'hb9df: y = 16'hfe00;
			16'hb9e0: y = 16'hfe00;
			16'hb9e1: y = 16'hfe00;
			16'hb9e2: y = 16'hfe00;
			16'hb9e3: y = 16'hfe00;
			16'hb9e4: y = 16'hfe00;
			16'hb9e5: y = 16'hfe00;
			16'hb9e6: y = 16'hfe00;
			16'hb9e7: y = 16'hfe00;
			16'hb9e8: y = 16'hfe00;
			16'hb9e9: y = 16'hfe00;
			16'hb9ea: y = 16'hfe00;
			16'hb9eb: y = 16'hfe00;
			16'hb9ec: y = 16'hfe00;
			16'hb9ed: y = 16'hfe00;
			16'hb9ee: y = 16'hfe00;
			16'hb9ef: y = 16'hfe00;
			16'hb9f0: y = 16'hfe00;
			16'hb9f1: y = 16'hfe00;
			16'hb9f2: y = 16'hfe00;
			16'hb9f3: y = 16'hfe00;
			16'hb9f4: y = 16'hfe00;
			16'hb9f5: y = 16'hfe00;
			16'hb9f6: y = 16'hfe00;
			16'hb9f7: y = 16'hfe00;
			16'hb9f8: y = 16'hfe00;
			16'hb9f9: y = 16'hfe00;
			16'hb9fa: y = 16'hfe00;
			16'hb9fb: y = 16'hfe00;
			16'hb9fc: y = 16'hfe00;
			16'hb9fd: y = 16'hfe00;
			16'hb9fe: y = 16'hfe00;
			16'hb9ff: y = 16'hfe00;
			16'hba00: y = 16'hfe00;
			16'hba01: y = 16'hfe00;
			16'hba02: y = 16'hfe00;
			16'hba03: y = 16'hfe00;
			16'hba04: y = 16'hfe00;
			16'hba05: y = 16'hfe00;
			16'hba06: y = 16'hfe00;
			16'hba07: y = 16'hfe00;
			16'hba08: y = 16'hfe00;
			16'hba09: y = 16'hfe00;
			16'hba0a: y = 16'hfe00;
			16'hba0b: y = 16'hfe00;
			16'hba0c: y = 16'hfe00;
			16'hba0d: y = 16'hfe00;
			16'hba0e: y = 16'hfe00;
			16'hba0f: y = 16'hfe00;
			16'hba10: y = 16'hfe00;
			16'hba11: y = 16'hfe00;
			16'hba12: y = 16'hfe00;
			16'hba13: y = 16'hfe00;
			16'hba14: y = 16'hfe00;
			16'hba15: y = 16'hfe00;
			16'hba16: y = 16'hfe00;
			16'hba17: y = 16'hfe00;
			16'hba18: y = 16'hfe00;
			16'hba19: y = 16'hfe00;
			16'hba1a: y = 16'hfe00;
			16'hba1b: y = 16'hfe00;
			16'hba1c: y = 16'hfe00;
			16'hba1d: y = 16'hfe00;
			16'hba1e: y = 16'hfe00;
			16'hba1f: y = 16'hfe00;
			16'hba20: y = 16'hfe00;
			16'hba21: y = 16'hfe00;
			16'hba22: y = 16'hfe00;
			16'hba23: y = 16'hfe00;
			16'hba24: y = 16'hfe00;
			16'hba25: y = 16'hfe00;
			16'hba26: y = 16'hfe00;
			16'hba27: y = 16'hfe00;
			16'hba28: y = 16'hfe00;
			16'hba29: y = 16'hfe00;
			16'hba2a: y = 16'hfe00;
			16'hba2b: y = 16'hfe00;
			16'hba2c: y = 16'hfe00;
			16'hba2d: y = 16'hfe00;
			16'hba2e: y = 16'hfe00;
			16'hba2f: y = 16'hfe00;
			16'hba30: y = 16'hfe00;
			16'hba31: y = 16'hfe00;
			16'hba32: y = 16'hfe00;
			16'hba33: y = 16'hfe00;
			16'hba34: y = 16'hfe00;
			16'hba35: y = 16'hfe00;
			16'hba36: y = 16'hfe00;
			16'hba37: y = 16'hfe00;
			16'hba38: y = 16'hfe00;
			16'hba39: y = 16'hfe00;
			16'hba3a: y = 16'hfe00;
			16'hba3b: y = 16'hfe00;
			16'hba3c: y = 16'hfe00;
			16'hba3d: y = 16'hfe00;
			16'hba3e: y = 16'hfe00;
			16'hba3f: y = 16'hfe00;
			16'hba40: y = 16'hfe00;
			16'hba41: y = 16'hfe00;
			16'hba42: y = 16'hfe00;
			16'hba43: y = 16'hfe00;
			16'hba44: y = 16'hfe00;
			16'hba45: y = 16'hfe00;
			16'hba46: y = 16'hfe00;
			16'hba47: y = 16'hfe00;
			16'hba48: y = 16'hfe00;
			16'hba49: y = 16'hfe00;
			16'hba4a: y = 16'hfe00;
			16'hba4b: y = 16'hfe00;
			16'hba4c: y = 16'hfe00;
			16'hba4d: y = 16'hfe00;
			16'hba4e: y = 16'hfe00;
			16'hba4f: y = 16'hfe00;
			16'hba50: y = 16'hfe00;
			16'hba51: y = 16'hfe00;
			16'hba52: y = 16'hfe00;
			16'hba53: y = 16'hfe00;
			16'hba54: y = 16'hfe00;
			16'hba55: y = 16'hfe00;
			16'hba56: y = 16'hfe00;
			16'hba57: y = 16'hfe00;
			16'hba58: y = 16'hfe00;
			16'hba59: y = 16'hfe00;
			16'hba5a: y = 16'hfe00;
			16'hba5b: y = 16'hfe00;
			16'hba5c: y = 16'hfe00;
			16'hba5d: y = 16'hfe00;
			16'hba5e: y = 16'hfe00;
			16'hba5f: y = 16'hfe00;
			16'hba60: y = 16'hfe00;
			16'hba61: y = 16'hfe00;
			16'hba62: y = 16'hfe00;
			16'hba63: y = 16'hfe00;
			16'hba64: y = 16'hfe00;
			16'hba65: y = 16'hfe00;
			16'hba66: y = 16'hfe00;
			16'hba67: y = 16'hfe00;
			16'hba68: y = 16'hfe00;
			16'hba69: y = 16'hfe00;
			16'hba6a: y = 16'hfe00;
			16'hba6b: y = 16'hfe00;
			16'hba6c: y = 16'hfe00;
			16'hba6d: y = 16'hfe00;
			16'hba6e: y = 16'hfe00;
			16'hba6f: y = 16'hfe00;
			16'hba70: y = 16'hfe00;
			16'hba71: y = 16'hfe00;
			16'hba72: y = 16'hfe00;
			16'hba73: y = 16'hfe00;
			16'hba74: y = 16'hfe00;
			16'hba75: y = 16'hfe00;
			16'hba76: y = 16'hfe00;
			16'hba77: y = 16'hfe00;
			16'hba78: y = 16'hfe00;
			16'hba79: y = 16'hfe00;
			16'hba7a: y = 16'hfe00;
			16'hba7b: y = 16'hfe00;
			16'hba7c: y = 16'hfe00;
			16'hba7d: y = 16'hfe00;
			16'hba7e: y = 16'hfe00;
			16'hba7f: y = 16'hfe00;
			16'hba80: y = 16'hfe00;
			16'hba81: y = 16'hfe00;
			16'hba82: y = 16'hfe00;
			16'hba83: y = 16'hfe00;
			16'hba84: y = 16'hfe00;
			16'hba85: y = 16'hfe00;
			16'hba86: y = 16'hfe00;
			16'hba87: y = 16'hfe00;
			16'hba88: y = 16'hfe00;
			16'hba89: y = 16'hfe00;
			16'hba8a: y = 16'hfe00;
			16'hba8b: y = 16'hfe00;
			16'hba8c: y = 16'hfe00;
			16'hba8d: y = 16'hfe00;
			16'hba8e: y = 16'hfe00;
			16'hba8f: y = 16'hfe00;
			16'hba90: y = 16'hfe00;
			16'hba91: y = 16'hfe00;
			16'hba92: y = 16'hfe00;
			16'hba93: y = 16'hfe00;
			16'hba94: y = 16'hfe00;
			16'hba95: y = 16'hfe00;
			16'hba96: y = 16'hfe00;
			16'hba97: y = 16'hfe00;
			16'hba98: y = 16'hfe00;
			16'hba99: y = 16'hfe00;
			16'hba9a: y = 16'hfe00;
			16'hba9b: y = 16'hfe00;
			16'hba9c: y = 16'hfe00;
			16'hba9d: y = 16'hfe00;
			16'hba9e: y = 16'hfe00;
			16'hba9f: y = 16'hfe00;
			16'hbaa0: y = 16'hfe00;
			16'hbaa1: y = 16'hfe00;
			16'hbaa2: y = 16'hfe00;
			16'hbaa3: y = 16'hfe00;
			16'hbaa4: y = 16'hfe00;
			16'hbaa5: y = 16'hfe00;
			16'hbaa6: y = 16'hfe00;
			16'hbaa7: y = 16'hfe00;
			16'hbaa8: y = 16'hfe00;
			16'hbaa9: y = 16'hfe00;
			16'hbaaa: y = 16'hfe00;
			16'hbaab: y = 16'hfe00;
			16'hbaac: y = 16'hfe00;
			16'hbaad: y = 16'hfe00;
			16'hbaae: y = 16'hfe00;
			16'hbaaf: y = 16'hfe00;
			16'hbab0: y = 16'hfe00;
			16'hbab1: y = 16'hfe00;
			16'hbab2: y = 16'hfe00;
			16'hbab3: y = 16'hfe00;
			16'hbab4: y = 16'hfe00;
			16'hbab5: y = 16'hfe00;
			16'hbab6: y = 16'hfe00;
			16'hbab7: y = 16'hfe00;
			16'hbab8: y = 16'hfe00;
			16'hbab9: y = 16'hfe00;
			16'hbaba: y = 16'hfe00;
			16'hbabb: y = 16'hfe00;
			16'hbabc: y = 16'hfe00;
			16'hbabd: y = 16'hfe00;
			16'hbabe: y = 16'hfe00;
			16'hbabf: y = 16'hfe00;
			16'hbac0: y = 16'hfe00;
			16'hbac1: y = 16'hfe00;
			16'hbac2: y = 16'hfe00;
			16'hbac3: y = 16'hfe00;
			16'hbac4: y = 16'hfe00;
			16'hbac5: y = 16'hfe00;
			16'hbac6: y = 16'hfe00;
			16'hbac7: y = 16'hfe00;
			16'hbac8: y = 16'hfe00;
			16'hbac9: y = 16'hfe00;
			16'hbaca: y = 16'hfe00;
			16'hbacb: y = 16'hfe00;
			16'hbacc: y = 16'hfe00;
			16'hbacd: y = 16'hfe00;
			16'hbace: y = 16'hfe00;
			16'hbacf: y = 16'hfe00;
			16'hbad0: y = 16'hfe00;
			16'hbad1: y = 16'hfe00;
			16'hbad2: y = 16'hfe00;
			16'hbad3: y = 16'hfe00;
			16'hbad4: y = 16'hfe00;
			16'hbad5: y = 16'hfe00;
			16'hbad6: y = 16'hfe00;
			16'hbad7: y = 16'hfe00;
			16'hbad8: y = 16'hfe00;
			16'hbad9: y = 16'hfe00;
			16'hbada: y = 16'hfe00;
			16'hbadb: y = 16'hfe00;
			16'hbadc: y = 16'hfe00;
			16'hbadd: y = 16'hfe00;
			16'hbade: y = 16'hfe00;
			16'hbadf: y = 16'hfe00;
			16'hbae0: y = 16'hfe00;
			16'hbae1: y = 16'hfe00;
			16'hbae2: y = 16'hfe00;
			16'hbae3: y = 16'hfe00;
			16'hbae4: y = 16'hfe00;
			16'hbae5: y = 16'hfe00;
			16'hbae6: y = 16'hfe00;
			16'hbae7: y = 16'hfe00;
			16'hbae8: y = 16'hfe00;
			16'hbae9: y = 16'hfe00;
			16'hbaea: y = 16'hfe00;
			16'hbaeb: y = 16'hfe00;
			16'hbaec: y = 16'hfe00;
			16'hbaed: y = 16'hfe00;
			16'hbaee: y = 16'hfe00;
			16'hbaef: y = 16'hfe00;
			16'hbaf0: y = 16'hfe00;
			16'hbaf1: y = 16'hfe00;
			16'hbaf2: y = 16'hfe00;
			16'hbaf3: y = 16'hfe00;
			16'hbaf4: y = 16'hfe00;
			16'hbaf5: y = 16'hfe00;
			16'hbaf6: y = 16'hfe00;
			16'hbaf7: y = 16'hfe00;
			16'hbaf8: y = 16'hfe00;
			16'hbaf9: y = 16'hfe00;
			16'hbafa: y = 16'hfe00;
			16'hbafb: y = 16'hfe00;
			16'hbafc: y = 16'hfe00;
			16'hbafd: y = 16'hfe00;
			16'hbafe: y = 16'hfe00;
			16'hbaff: y = 16'hfe00;
			16'hbb00: y = 16'hfe00;
			16'hbb01: y = 16'hfe00;
			16'hbb02: y = 16'hfe00;
			16'hbb03: y = 16'hfe00;
			16'hbb04: y = 16'hfe00;
			16'hbb05: y = 16'hfe00;
			16'hbb06: y = 16'hfe00;
			16'hbb07: y = 16'hfe00;
			16'hbb08: y = 16'hfe00;
			16'hbb09: y = 16'hfe00;
			16'hbb0a: y = 16'hfe00;
			16'hbb0b: y = 16'hfe00;
			16'hbb0c: y = 16'hfe00;
			16'hbb0d: y = 16'hfe00;
			16'hbb0e: y = 16'hfe00;
			16'hbb0f: y = 16'hfe00;
			16'hbb10: y = 16'hfe00;
			16'hbb11: y = 16'hfe00;
			16'hbb12: y = 16'hfe00;
			16'hbb13: y = 16'hfe00;
			16'hbb14: y = 16'hfe00;
			16'hbb15: y = 16'hfe00;
			16'hbb16: y = 16'hfe00;
			16'hbb17: y = 16'hfe00;
			16'hbb18: y = 16'hfe00;
			16'hbb19: y = 16'hfe00;
			16'hbb1a: y = 16'hfe00;
			16'hbb1b: y = 16'hfe00;
			16'hbb1c: y = 16'hfe00;
			16'hbb1d: y = 16'hfe00;
			16'hbb1e: y = 16'hfe00;
			16'hbb1f: y = 16'hfe00;
			16'hbb20: y = 16'hfe00;
			16'hbb21: y = 16'hfe00;
			16'hbb22: y = 16'hfe00;
			16'hbb23: y = 16'hfe00;
			16'hbb24: y = 16'hfe00;
			16'hbb25: y = 16'hfe00;
			16'hbb26: y = 16'hfe00;
			16'hbb27: y = 16'hfe00;
			16'hbb28: y = 16'hfe00;
			16'hbb29: y = 16'hfe00;
			16'hbb2a: y = 16'hfe00;
			16'hbb2b: y = 16'hfe00;
			16'hbb2c: y = 16'hfe00;
			16'hbb2d: y = 16'hfe00;
			16'hbb2e: y = 16'hfe00;
			16'hbb2f: y = 16'hfe00;
			16'hbb30: y = 16'hfe00;
			16'hbb31: y = 16'hfe00;
			16'hbb32: y = 16'hfe00;
			16'hbb33: y = 16'hfe00;
			16'hbb34: y = 16'hfe00;
			16'hbb35: y = 16'hfe00;
			16'hbb36: y = 16'hfe00;
			16'hbb37: y = 16'hfe00;
			16'hbb38: y = 16'hfe00;
			16'hbb39: y = 16'hfe00;
			16'hbb3a: y = 16'hfe00;
			16'hbb3b: y = 16'hfe00;
			16'hbb3c: y = 16'hfe00;
			16'hbb3d: y = 16'hfe00;
			16'hbb3e: y = 16'hfe00;
			16'hbb3f: y = 16'hfe00;
			16'hbb40: y = 16'hfe00;
			16'hbb41: y = 16'hfe00;
			16'hbb42: y = 16'hfe00;
			16'hbb43: y = 16'hfe00;
			16'hbb44: y = 16'hfe00;
			16'hbb45: y = 16'hfe00;
			16'hbb46: y = 16'hfe00;
			16'hbb47: y = 16'hfe00;
			16'hbb48: y = 16'hfe00;
			16'hbb49: y = 16'hfe00;
			16'hbb4a: y = 16'hfe00;
			16'hbb4b: y = 16'hfe00;
			16'hbb4c: y = 16'hfe00;
			16'hbb4d: y = 16'hfe00;
			16'hbb4e: y = 16'hfe00;
			16'hbb4f: y = 16'hfe00;
			16'hbb50: y = 16'hfe00;
			16'hbb51: y = 16'hfe00;
			16'hbb52: y = 16'hfe00;
			16'hbb53: y = 16'hfe00;
			16'hbb54: y = 16'hfe00;
			16'hbb55: y = 16'hfe00;
			16'hbb56: y = 16'hfe00;
			16'hbb57: y = 16'hfe00;
			16'hbb58: y = 16'hfe00;
			16'hbb59: y = 16'hfe00;
			16'hbb5a: y = 16'hfe00;
			16'hbb5b: y = 16'hfe00;
			16'hbb5c: y = 16'hfe00;
			16'hbb5d: y = 16'hfe00;
			16'hbb5e: y = 16'hfe00;
			16'hbb5f: y = 16'hfe00;
			16'hbb60: y = 16'hfe00;
			16'hbb61: y = 16'hfe00;
			16'hbb62: y = 16'hfe00;
			16'hbb63: y = 16'hfe00;
			16'hbb64: y = 16'hfe00;
			16'hbb65: y = 16'hfe00;
			16'hbb66: y = 16'hfe00;
			16'hbb67: y = 16'hfe00;
			16'hbb68: y = 16'hfe00;
			16'hbb69: y = 16'hfe00;
			16'hbb6a: y = 16'hfe00;
			16'hbb6b: y = 16'hfe00;
			16'hbb6c: y = 16'hfe00;
			16'hbb6d: y = 16'hfe00;
			16'hbb6e: y = 16'hfe00;
			16'hbb6f: y = 16'hfe00;
			16'hbb70: y = 16'hfe00;
			16'hbb71: y = 16'hfe00;
			16'hbb72: y = 16'hfe00;
			16'hbb73: y = 16'hfe00;
			16'hbb74: y = 16'hfe00;
			16'hbb75: y = 16'hfe00;
			16'hbb76: y = 16'hfe00;
			16'hbb77: y = 16'hfe00;
			16'hbb78: y = 16'hfe00;
			16'hbb79: y = 16'hfe00;
			16'hbb7a: y = 16'hfe00;
			16'hbb7b: y = 16'hfe00;
			16'hbb7c: y = 16'hfe00;
			16'hbb7d: y = 16'hfe00;
			16'hbb7e: y = 16'hfe00;
			16'hbb7f: y = 16'hfe00;
			16'hbb80: y = 16'hfe00;
			16'hbb81: y = 16'hfe00;
			16'hbb82: y = 16'hfe00;
			16'hbb83: y = 16'hfe00;
			16'hbb84: y = 16'hfe00;
			16'hbb85: y = 16'hfe00;
			16'hbb86: y = 16'hfe00;
			16'hbb87: y = 16'hfe00;
			16'hbb88: y = 16'hfe00;
			16'hbb89: y = 16'hfe00;
			16'hbb8a: y = 16'hfe00;
			16'hbb8b: y = 16'hfe00;
			16'hbb8c: y = 16'hfe00;
			16'hbb8d: y = 16'hfe00;
			16'hbb8e: y = 16'hfe00;
			16'hbb8f: y = 16'hfe00;
			16'hbb90: y = 16'hfe00;
			16'hbb91: y = 16'hfe00;
			16'hbb92: y = 16'hfe00;
			16'hbb93: y = 16'hfe00;
			16'hbb94: y = 16'hfe00;
			16'hbb95: y = 16'hfe00;
			16'hbb96: y = 16'hfe00;
			16'hbb97: y = 16'hfe00;
			16'hbb98: y = 16'hfe00;
			16'hbb99: y = 16'hfe00;
			16'hbb9a: y = 16'hfe00;
			16'hbb9b: y = 16'hfe00;
			16'hbb9c: y = 16'hfe00;
			16'hbb9d: y = 16'hfe00;
			16'hbb9e: y = 16'hfe00;
			16'hbb9f: y = 16'hfe00;
			16'hbba0: y = 16'hfe00;
			16'hbba1: y = 16'hfe00;
			16'hbba2: y = 16'hfe00;
			16'hbba3: y = 16'hfe00;
			16'hbba4: y = 16'hfe00;
			16'hbba5: y = 16'hfe00;
			16'hbba6: y = 16'hfe00;
			16'hbba7: y = 16'hfe00;
			16'hbba8: y = 16'hfe00;
			16'hbba9: y = 16'hfe00;
			16'hbbaa: y = 16'hfe00;
			16'hbbab: y = 16'hfe00;
			16'hbbac: y = 16'hfe00;
			16'hbbad: y = 16'hfe00;
			16'hbbae: y = 16'hfe00;
			16'hbbaf: y = 16'hfe00;
			16'hbbb0: y = 16'hfe00;
			16'hbbb1: y = 16'hfe00;
			16'hbbb2: y = 16'hfe00;
			16'hbbb3: y = 16'hfe00;
			16'hbbb4: y = 16'hfe00;
			16'hbbb5: y = 16'hfe00;
			16'hbbb6: y = 16'hfe00;
			16'hbbb7: y = 16'hfe00;
			16'hbbb8: y = 16'hfe00;
			16'hbbb9: y = 16'hfe00;
			16'hbbba: y = 16'hfe00;
			16'hbbbb: y = 16'hfe00;
			16'hbbbc: y = 16'hfe00;
			16'hbbbd: y = 16'hfe00;
			16'hbbbe: y = 16'hfe00;
			16'hbbbf: y = 16'hfe00;
			16'hbbc0: y = 16'hfe00;
			16'hbbc1: y = 16'hfe00;
			16'hbbc2: y = 16'hfe00;
			16'hbbc3: y = 16'hfe00;
			16'hbbc4: y = 16'hfe00;
			16'hbbc5: y = 16'hfe00;
			16'hbbc6: y = 16'hfe00;
			16'hbbc7: y = 16'hfe00;
			16'hbbc8: y = 16'hfe00;
			16'hbbc9: y = 16'hfe00;
			16'hbbca: y = 16'hfe00;
			16'hbbcb: y = 16'hfe00;
			16'hbbcc: y = 16'hfe00;
			16'hbbcd: y = 16'hfe00;
			16'hbbce: y = 16'hfe00;
			16'hbbcf: y = 16'hfe00;
			16'hbbd0: y = 16'hfe00;
			16'hbbd1: y = 16'hfe00;
			16'hbbd2: y = 16'hfe00;
			16'hbbd3: y = 16'hfe00;
			16'hbbd4: y = 16'hfe00;
			16'hbbd5: y = 16'hfe00;
			16'hbbd6: y = 16'hfe00;
			16'hbbd7: y = 16'hfe00;
			16'hbbd8: y = 16'hfe00;
			16'hbbd9: y = 16'hfe00;
			16'hbbda: y = 16'hfe00;
			16'hbbdb: y = 16'hfe00;
			16'hbbdc: y = 16'hfe00;
			16'hbbdd: y = 16'hfe00;
			16'hbbde: y = 16'hfe00;
			16'hbbdf: y = 16'hfe00;
			16'hbbe0: y = 16'hfe00;
			16'hbbe1: y = 16'hfe00;
			16'hbbe2: y = 16'hfe00;
			16'hbbe3: y = 16'hfe00;
			16'hbbe4: y = 16'hfe00;
			16'hbbe5: y = 16'hfe00;
			16'hbbe6: y = 16'hfe00;
			16'hbbe7: y = 16'hfe00;
			16'hbbe8: y = 16'hfe00;
			16'hbbe9: y = 16'hfe00;
			16'hbbea: y = 16'hfe00;
			16'hbbeb: y = 16'hfe00;
			16'hbbec: y = 16'hfe00;
			16'hbbed: y = 16'hfe00;
			16'hbbee: y = 16'hfe00;
			16'hbbef: y = 16'hfe00;
			16'hbbf0: y = 16'hfe00;
			16'hbbf1: y = 16'hfe00;
			16'hbbf2: y = 16'hfe00;
			16'hbbf3: y = 16'hfe00;
			16'hbbf4: y = 16'hfe00;
			16'hbbf5: y = 16'hfe00;
			16'hbbf6: y = 16'hfe00;
			16'hbbf7: y = 16'hfe00;
			16'hbbf8: y = 16'hfe00;
			16'hbbf9: y = 16'hfe00;
			16'hbbfa: y = 16'hfe00;
			16'hbbfb: y = 16'hfe00;
			16'hbbfc: y = 16'hfe00;
			16'hbbfd: y = 16'hfe00;
			16'hbbfe: y = 16'hfe00;
			16'hbbff: y = 16'hfe00;
			16'hbc00: y = 16'hfe00;
			16'hbc01: y = 16'hfe00;
			16'hbc02: y = 16'hfe00;
			16'hbc03: y = 16'hfe00;
			16'hbc04: y = 16'hfe00;
			16'hbc05: y = 16'hfe00;
			16'hbc06: y = 16'hfe00;
			16'hbc07: y = 16'hfe00;
			16'hbc08: y = 16'hfe00;
			16'hbc09: y = 16'hfe00;
			16'hbc0a: y = 16'hfe00;
			16'hbc0b: y = 16'hfe00;
			16'hbc0c: y = 16'hfe00;
			16'hbc0d: y = 16'hfe00;
			16'hbc0e: y = 16'hfe00;
			16'hbc0f: y = 16'hfe00;
			16'hbc10: y = 16'hfe00;
			16'hbc11: y = 16'hfe00;
			16'hbc12: y = 16'hfe00;
			16'hbc13: y = 16'hfe00;
			16'hbc14: y = 16'hfe00;
			16'hbc15: y = 16'hfe00;
			16'hbc16: y = 16'hfe00;
			16'hbc17: y = 16'hfe00;
			16'hbc18: y = 16'hfe00;
			16'hbc19: y = 16'hfe00;
			16'hbc1a: y = 16'hfe00;
			16'hbc1b: y = 16'hfe00;
			16'hbc1c: y = 16'hfe00;
			16'hbc1d: y = 16'hfe00;
			16'hbc1e: y = 16'hfe00;
			16'hbc1f: y = 16'hfe00;
			16'hbc20: y = 16'hfe00;
			16'hbc21: y = 16'hfe00;
			16'hbc22: y = 16'hfe00;
			16'hbc23: y = 16'hfe00;
			16'hbc24: y = 16'hfe00;
			16'hbc25: y = 16'hfe00;
			16'hbc26: y = 16'hfe00;
			16'hbc27: y = 16'hfe00;
			16'hbc28: y = 16'hfe00;
			16'hbc29: y = 16'hfe00;
			16'hbc2a: y = 16'hfe00;
			16'hbc2b: y = 16'hfe00;
			16'hbc2c: y = 16'hfe00;
			16'hbc2d: y = 16'hfe00;
			16'hbc2e: y = 16'hfe00;
			16'hbc2f: y = 16'hfe00;
			16'hbc30: y = 16'hfe00;
			16'hbc31: y = 16'hfe00;
			16'hbc32: y = 16'hfe00;
			16'hbc33: y = 16'hfe00;
			16'hbc34: y = 16'hfe00;
			16'hbc35: y = 16'hfe00;
			16'hbc36: y = 16'hfe00;
			16'hbc37: y = 16'hfe00;
			16'hbc38: y = 16'hfe00;
			16'hbc39: y = 16'hfe00;
			16'hbc3a: y = 16'hfe00;
			16'hbc3b: y = 16'hfe00;
			16'hbc3c: y = 16'hfe00;
			16'hbc3d: y = 16'hfe00;
			16'hbc3e: y = 16'hfe00;
			16'hbc3f: y = 16'hfe00;
			16'hbc40: y = 16'hfe00;
			16'hbc41: y = 16'hfe00;
			16'hbc42: y = 16'hfe00;
			16'hbc43: y = 16'hfe00;
			16'hbc44: y = 16'hfe00;
			16'hbc45: y = 16'hfe00;
			16'hbc46: y = 16'hfe00;
			16'hbc47: y = 16'hfe00;
			16'hbc48: y = 16'hfe00;
			16'hbc49: y = 16'hfe00;
			16'hbc4a: y = 16'hfe00;
			16'hbc4b: y = 16'hfe00;
			16'hbc4c: y = 16'hfe00;
			16'hbc4d: y = 16'hfe00;
			16'hbc4e: y = 16'hfe00;
			16'hbc4f: y = 16'hfe00;
			16'hbc50: y = 16'hfe00;
			16'hbc51: y = 16'hfe00;
			16'hbc52: y = 16'hfe00;
			16'hbc53: y = 16'hfe00;
			16'hbc54: y = 16'hfe00;
			16'hbc55: y = 16'hfe00;
			16'hbc56: y = 16'hfe00;
			16'hbc57: y = 16'hfe00;
			16'hbc58: y = 16'hfe00;
			16'hbc59: y = 16'hfe00;
			16'hbc5a: y = 16'hfe00;
			16'hbc5b: y = 16'hfe00;
			16'hbc5c: y = 16'hfe00;
			16'hbc5d: y = 16'hfe00;
			16'hbc5e: y = 16'hfe00;
			16'hbc5f: y = 16'hfe00;
			16'hbc60: y = 16'hfe00;
			16'hbc61: y = 16'hfe00;
			16'hbc62: y = 16'hfe00;
			16'hbc63: y = 16'hfe00;
			16'hbc64: y = 16'hfe00;
			16'hbc65: y = 16'hfe00;
			16'hbc66: y = 16'hfe00;
			16'hbc67: y = 16'hfe00;
			16'hbc68: y = 16'hfe00;
			16'hbc69: y = 16'hfe00;
			16'hbc6a: y = 16'hfe00;
			16'hbc6b: y = 16'hfe00;
			16'hbc6c: y = 16'hfe00;
			16'hbc6d: y = 16'hfe00;
			16'hbc6e: y = 16'hfe00;
			16'hbc6f: y = 16'hfe00;
			16'hbc70: y = 16'hfe00;
			16'hbc71: y = 16'hfe00;
			16'hbc72: y = 16'hfe00;
			16'hbc73: y = 16'hfe00;
			16'hbc74: y = 16'hfe00;
			16'hbc75: y = 16'hfe00;
			16'hbc76: y = 16'hfe00;
			16'hbc77: y = 16'hfe00;
			16'hbc78: y = 16'hfe00;
			16'hbc79: y = 16'hfe00;
			16'hbc7a: y = 16'hfe00;
			16'hbc7b: y = 16'hfe00;
			16'hbc7c: y = 16'hfe00;
			16'hbc7d: y = 16'hfe00;
			16'hbc7e: y = 16'hfe00;
			16'hbc7f: y = 16'hfe00;
			16'hbc80: y = 16'hfe00;
			16'hbc81: y = 16'hfe00;
			16'hbc82: y = 16'hfe00;
			16'hbc83: y = 16'hfe00;
			16'hbc84: y = 16'hfe00;
			16'hbc85: y = 16'hfe00;
			16'hbc86: y = 16'hfe00;
			16'hbc87: y = 16'hfe00;
			16'hbc88: y = 16'hfe00;
			16'hbc89: y = 16'hfe00;
			16'hbc8a: y = 16'hfe00;
			16'hbc8b: y = 16'hfe00;
			16'hbc8c: y = 16'hfe00;
			16'hbc8d: y = 16'hfe00;
			16'hbc8e: y = 16'hfe00;
			16'hbc8f: y = 16'hfe00;
			16'hbc90: y = 16'hfe00;
			16'hbc91: y = 16'hfe00;
			16'hbc92: y = 16'hfe00;
			16'hbc93: y = 16'hfe00;
			16'hbc94: y = 16'hfe00;
			16'hbc95: y = 16'hfe00;
			16'hbc96: y = 16'hfe00;
			16'hbc97: y = 16'hfe00;
			16'hbc98: y = 16'hfe00;
			16'hbc99: y = 16'hfe00;
			16'hbc9a: y = 16'hfe00;
			16'hbc9b: y = 16'hfe00;
			16'hbc9c: y = 16'hfe00;
			16'hbc9d: y = 16'hfe00;
			16'hbc9e: y = 16'hfe00;
			16'hbc9f: y = 16'hfe00;
			16'hbca0: y = 16'hfe00;
			16'hbca1: y = 16'hfe00;
			16'hbca2: y = 16'hfe00;
			16'hbca3: y = 16'hfe00;
			16'hbca4: y = 16'hfe00;
			16'hbca5: y = 16'hfe00;
			16'hbca6: y = 16'hfe00;
			16'hbca7: y = 16'hfe00;
			16'hbca8: y = 16'hfe00;
			16'hbca9: y = 16'hfe00;
			16'hbcaa: y = 16'hfe00;
			16'hbcab: y = 16'hfe00;
			16'hbcac: y = 16'hfe00;
			16'hbcad: y = 16'hfe00;
			16'hbcae: y = 16'hfe00;
			16'hbcaf: y = 16'hfe00;
			16'hbcb0: y = 16'hfe00;
			16'hbcb1: y = 16'hfe00;
			16'hbcb2: y = 16'hfe00;
			16'hbcb3: y = 16'hfe00;
			16'hbcb4: y = 16'hfe00;
			16'hbcb5: y = 16'hfe00;
			16'hbcb6: y = 16'hfe00;
			16'hbcb7: y = 16'hfe00;
			16'hbcb8: y = 16'hfe00;
			16'hbcb9: y = 16'hfe00;
			16'hbcba: y = 16'hfe00;
			16'hbcbb: y = 16'hfe00;
			16'hbcbc: y = 16'hfe00;
			16'hbcbd: y = 16'hfe00;
			16'hbcbe: y = 16'hfe00;
			16'hbcbf: y = 16'hfe00;
			16'hbcc0: y = 16'hfe00;
			16'hbcc1: y = 16'hfe00;
			16'hbcc2: y = 16'hfe00;
			16'hbcc3: y = 16'hfe00;
			16'hbcc4: y = 16'hfe00;
			16'hbcc5: y = 16'hfe00;
			16'hbcc6: y = 16'hfe00;
			16'hbcc7: y = 16'hfe00;
			16'hbcc8: y = 16'hfe00;
			16'hbcc9: y = 16'hfe00;
			16'hbcca: y = 16'hfe00;
			16'hbccb: y = 16'hfe00;
			16'hbccc: y = 16'hfe00;
			16'hbccd: y = 16'hfe00;
			16'hbcce: y = 16'hfe00;
			16'hbccf: y = 16'hfe00;
			16'hbcd0: y = 16'hfe00;
			16'hbcd1: y = 16'hfe00;
			16'hbcd2: y = 16'hfe00;
			16'hbcd3: y = 16'hfe00;
			16'hbcd4: y = 16'hfe00;
			16'hbcd5: y = 16'hfe00;
			16'hbcd6: y = 16'hfe00;
			16'hbcd7: y = 16'hfe00;
			16'hbcd8: y = 16'hfe00;
			16'hbcd9: y = 16'hfe00;
			16'hbcda: y = 16'hfe00;
			16'hbcdb: y = 16'hfe00;
			16'hbcdc: y = 16'hfe00;
			16'hbcdd: y = 16'hfe00;
			16'hbcde: y = 16'hfe00;
			16'hbcdf: y = 16'hfe00;
			16'hbce0: y = 16'hfe00;
			16'hbce1: y = 16'hfe00;
			16'hbce2: y = 16'hfe00;
			16'hbce3: y = 16'hfe00;
			16'hbce4: y = 16'hfe00;
			16'hbce5: y = 16'hfe00;
			16'hbce6: y = 16'hfe00;
			16'hbce7: y = 16'hfe00;
			16'hbce8: y = 16'hfe00;
			16'hbce9: y = 16'hfe00;
			16'hbcea: y = 16'hfe00;
			16'hbceb: y = 16'hfe00;
			16'hbcec: y = 16'hfe00;
			16'hbced: y = 16'hfe00;
			16'hbcee: y = 16'hfe00;
			16'hbcef: y = 16'hfe00;
			16'hbcf0: y = 16'hfe00;
			16'hbcf1: y = 16'hfe00;
			16'hbcf2: y = 16'hfe00;
			16'hbcf3: y = 16'hfe00;
			16'hbcf4: y = 16'hfe00;
			16'hbcf5: y = 16'hfe00;
			16'hbcf6: y = 16'hfe00;
			16'hbcf7: y = 16'hfe00;
			16'hbcf8: y = 16'hfe00;
			16'hbcf9: y = 16'hfe00;
			16'hbcfa: y = 16'hfe00;
			16'hbcfb: y = 16'hfe00;
			16'hbcfc: y = 16'hfe00;
			16'hbcfd: y = 16'hfe00;
			16'hbcfe: y = 16'hfe00;
			16'hbcff: y = 16'hfe00;
			16'hbd00: y = 16'hfe00;
			16'hbd01: y = 16'hfe00;
			16'hbd02: y = 16'hfe00;
			16'hbd03: y = 16'hfe00;
			16'hbd04: y = 16'hfe00;
			16'hbd05: y = 16'hfe00;
			16'hbd06: y = 16'hfe00;
			16'hbd07: y = 16'hfe00;
			16'hbd08: y = 16'hfe00;
			16'hbd09: y = 16'hfe00;
			16'hbd0a: y = 16'hfe00;
			16'hbd0b: y = 16'hfe00;
			16'hbd0c: y = 16'hfe00;
			16'hbd0d: y = 16'hfe00;
			16'hbd0e: y = 16'hfe00;
			16'hbd0f: y = 16'hfe00;
			16'hbd10: y = 16'hfe00;
			16'hbd11: y = 16'hfe00;
			16'hbd12: y = 16'hfe00;
			16'hbd13: y = 16'hfe00;
			16'hbd14: y = 16'hfe00;
			16'hbd15: y = 16'hfe00;
			16'hbd16: y = 16'hfe00;
			16'hbd17: y = 16'hfe00;
			16'hbd18: y = 16'hfe00;
			16'hbd19: y = 16'hfe00;
			16'hbd1a: y = 16'hfe00;
			16'hbd1b: y = 16'hfe00;
			16'hbd1c: y = 16'hfe00;
			16'hbd1d: y = 16'hfe00;
			16'hbd1e: y = 16'hfe00;
			16'hbd1f: y = 16'hfe00;
			16'hbd20: y = 16'hfe00;
			16'hbd21: y = 16'hfe00;
			16'hbd22: y = 16'hfe00;
			16'hbd23: y = 16'hfe00;
			16'hbd24: y = 16'hfe00;
			16'hbd25: y = 16'hfe00;
			16'hbd26: y = 16'hfe00;
			16'hbd27: y = 16'hfe00;
			16'hbd28: y = 16'hfe00;
			16'hbd29: y = 16'hfe00;
			16'hbd2a: y = 16'hfe00;
			16'hbd2b: y = 16'hfe00;
			16'hbd2c: y = 16'hfe00;
			16'hbd2d: y = 16'hfe00;
			16'hbd2e: y = 16'hfe00;
			16'hbd2f: y = 16'hfe00;
			16'hbd30: y = 16'hfe00;
			16'hbd31: y = 16'hfe00;
			16'hbd32: y = 16'hfe00;
			16'hbd33: y = 16'hfe00;
			16'hbd34: y = 16'hfe00;
			16'hbd35: y = 16'hfe00;
			16'hbd36: y = 16'hfe00;
			16'hbd37: y = 16'hfe00;
			16'hbd38: y = 16'hfe00;
			16'hbd39: y = 16'hfe00;
			16'hbd3a: y = 16'hfe00;
			16'hbd3b: y = 16'hfe00;
			16'hbd3c: y = 16'hfe00;
			16'hbd3d: y = 16'hfe00;
			16'hbd3e: y = 16'hfe00;
			16'hbd3f: y = 16'hfe00;
			16'hbd40: y = 16'hfe00;
			16'hbd41: y = 16'hfe00;
			16'hbd42: y = 16'hfe00;
			16'hbd43: y = 16'hfe00;
			16'hbd44: y = 16'hfe00;
			16'hbd45: y = 16'hfe00;
			16'hbd46: y = 16'hfe00;
			16'hbd47: y = 16'hfe00;
			16'hbd48: y = 16'hfe00;
			16'hbd49: y = 16'hfe00;
			16'hbd4a: y = 16'hfe00;
			16'hbd4b: y = 16'hfe00;
			16'hbd4c: y = 16'hfe00;
			16'hbd4d: y = 16'hfe00;
			16'hbd4e: y = 16'hfe00;
			16'hbd4f: y = 16'hfe00;
			16'hbd50: y = 16'hfe00;
			16'hbd51: y = 16'hfe00;
			16'hbd52: y = 16'hfe00;
			16'hbd53: y = 16'hfe00;
			16'hbd54: y = 16'hfe00;
			16'hbd55: y = 16'hfe00;
			16'hbd56: y = 16'hfe00;
			16'hbd57: y = 16'hfe00;
			16'hbd58: y = 16'hfe00;
			16'hbd59: y = 16'hfe00;
			16'hbd5a: y = 16'hfe00;
			16'hbd5b: y = 16'hfe00;
			16'hbd5c: y = 16'hfe00;
			16'hbd5d: y = 16'hfe00;
			16'hbd5e: y = 16'hfe00;
			16'hbd5f: y = 16'hfe00;
			16'hbd60: y = 16'hfe00;
			16'hbd61: y = 16'hfe00;
			16'hbd62: y = 16'hfe00;
			16'hbd63: y = 16'hfe00;
			16'hbd64: y = 16'hfe00;
			16'hbd65: y = 16'hfe00;
			16'hbd66: y = 16'hfe00;
			16'hbd67: y = 16'hfe00;
			16'hbd68: y = 16'hfe00;
			16'hbd69: y = 16'hfe00;
			16'hbd6a: y = 16'hfe00;
			16'hbd6b: y = 16'hfe00;
			16'hbd6c: y = 16'hfe00;
			16'hbd6d: y = 16'hfe00;
			16'hbd6e: y = 16'hfe00;
			16'hbd6f: y = 16'hfe00;
			16'hbd70: y = 16'hfe00;
			16'hbd71: y = 16'hfe00;
			16'hbd72: y = 16'hfe00;
			16'hbd73: y = 16'hfe00;
			16'hbd74: y = 16'hfe00;
			16'hbd75: y = 16'hfe00;
			16'hbd76: y = 16'hfe00;
			16'hbd77: y = 16'hfe00;
			16'hbd78: y = 16'hfe00;
			16'hbd79: y = 16'hfe00;
			16'hbd7a: y = 16'hfe00;
			16'hbd7b: y = 16'hfe00;
			16'hbd7c: y = 16'hfe00;
			16'hbd7d: y = 16'hfe00;
			16'hbd7e: y = 16'hfe00;
			16'hbd7f: y = 16'hfe00;
			16'hbd80: y = 16'hfe00;
			16'hbd81: y = 16'hfe00;
			16'hbd82: y = 16'hfe00;
			16'hbd83: y = 16'hfe00;
			16'hbd84: y = 16'hfe00;
			16'hbd85: y = 16'hfe00;
			16'hbd86: y = 16'hfe00;
			16'hbd87: y = 16'hfe00;
			16'hbd88: y = 16'hfe00;
			16'hbd89: y = 16'hfe00;
			16'hbd8a: y = 16'hfe00;
			16'hbd8b: y = 16'hfe00;
			16'hbd8c: y = 16'hfe00;
			16'hbd8d: y = 16'hfe00;
			16'hbd8e: y = 16'hfe00;
			16'hbd8f: y = 16'hfe00;
			16'hbd90: y = 16'hfe00;
			16'hbd91: y = 16'hfe00;
			16'hbd92: y = 16'hfe00;
			16'hbd93: y = 16'hfe00;
			16'hbd94: y = 16'hfe00;
			16'hbd95: y = 16'hfe00;
			16'hbd96: y = 16'hfe00;
			16'hbd97: y = 16'hfe00;
			16'hbd98: y = 16'hfe00;
			16'hbd99: y = 16'hfe00;
			16'hbd9a: y = 16'hfe00;
			16'hbd9b: y = 16'hfe00;
			16'hbd9c: y = 16'hfe00;
			16'hbd9d: y = 16'hfe00;
			16'hbd9e: y = 16'hfe00;
			16'hbd9f: y = 16'hfe00;
			16'hbda0: y = 16'hfe00;
			16'hbda1: y = 16'hfe00;
			16'hbda2: y = 16'hfe00;
			16'hbda3: y = 16'hfe00;
			16'hbda4: y = 16'hfe00;
			16'hbda5: y = 16'hfe00;
			16'hbda6: y = 16'hfe00;
			16'hbda7: y = 16'hfe00;
			16'hbda8: y = 16'hfe00;
			16'hbda9: y = 16'hfe00;
			16'hbdaa: y = 16'hfe00;
			16'hbdab: y = 16'hfe00;
			16'hbdac: y = 16'hfe00;
			16'hbdad: y = 16'hfe00;
			16'hbdae: y = 16'hfe00;
			16'hbdaf: y = 16'hfe00;
			16'hbdb0: y = 16'hfe00;
			16'hbdb1: y = 16'hfe00;
			16'hbdb2: y = 16'hfe00;
			16'hbdb3: y = 16'hfe00;
			16'hbdb4: y = 16'hfe00;
			16'hbdb5: y = 16'hfe00;
			16'hbdb6: y = 16'hfe00;
			16'hbdb7: y = 16'hfe00;
			16'hbdb8: y = 16'hfe00;
			16'hbdb9: y = 16'hfe00;
			16'hbdba: y = 16'hfe00;
			16'hbdbb: y = 16'hfe00;
			16'hbdbc: y = 16'hfe00;
			16'hbdbd: y = 16'hfe00;
			16'hbdbe: y = 16'hfe00;
			16'hbdbf: y = 16'hfe00;
			16'hbdc0: y = 16'hfe00;
			16'hbdc1: y = 16'hfe00;
			16'hbdc2: y = 16'hfe00;
			16'hbdc3: y = 16'hfe00;
			16'hbdc4: y = 16'hfe00;
			16'hbdc5: y = 16'hfe00;
			16'hbdc6: y = 16'hfe00;
			16'hbdc7: y = 16'hfe00;
			16'hbdc8: y = 16'hfe00;
			16'hbdc9: y = 16'hfe00;
			16'hbdca: y = 16'hfe00;
			16'hbdcb: y = 16'hfe00;
			16'hbdcc: y = 16'hfe00;
			16'hbdcd: y = 16'hfe00;
			16'hbdce: y = 16'hfe00;
			16'hbdcf: y = 16'hfe00;
			16'hbdd0: y = 16'hfe00;
			16'hbdd1: y = 16'hfe00;
			16'hbdd2: y = 16'hfe00;
			16'hbdd3: y = 16'hfe00;
			16'hbdd4: y = 16'hfe00;
			16'hbdd5: y = 16'hfe00;
			16'hbdd6: y = 16'hfe00;
			16'hbdd7: y = 16'hfe00;
			16'hbdd8: y = 16'hfe00;
			16'hbdd9: y = 16'hfe00;
			16'hbdda: y = 16'hfe00;
			16'hbddb: y = 16'hfe00;
			16'hbddc: y = 16'hfe00;
			16'hbddd: y = 16'hfe00;
			16'hbdde: y = 16'hfe00;
			16'hbddf: y = 16'hfe00;
			16'hbde0: y = 16'hfe00;
			16'hbde1: y = 16'hfe00;
			16'hbde2: y = 16'hfe00;
			16'hbde3: y = 16'hfe00;
			16'hbde4: y = 16'hfe00;
			16'hbde5: y = 16'hfe00;
			16'hbde6: y = 16'hfe00;
			16'hbde7: y = 16'hfe00;
			16'hbde8: y = 16'hfe00;
			16'hbde9: y = 16'hfe00;
			16'hbdea: y = 16'hfe00;
			16'hbdeb: y = 16'hfe00;
			16'hbdec: y = 16'hfe00;
			16'hbded: y = 16'hfe00;
			16'hbdee: y = 16'hfe00;
			16'hbdef: y = 16'hfe00;
			16'hbdf0: y = 16'hfe00;
			16'hbdf1: y = 16'hfe00;
			16'hbdf2: y = 16'hfe00;
			16'hbdf3: y = 16'hfe00;
			16'hbdf4: y = 16'hfe00;
			16'hbdf5: y = 16'hfe00;
			16'hbdf6: y = 16'hfe00;
			16'hbdf7: y = 16'hfe00;
			16'hbdf8: y = 16'hfe00;
			16'hbdf9: y = 16'hfe00;
			16'hbdfa: y = 16'hfe00;
			16'hbdfb: y = 16'hfe00;
			16'hbdfc: y = 16'hfe00;
			16'hbdfd: y = 16'hfe00;
			16'hbdfe: y = 16'hfe00;
			16'hbdff: y = 16'hfe00;
			16'hbe00: y = 16'hfe00;
			16'hbe01: y = 16'hfe00;
			16'hbe02: y = 16'hfe00;
			16'hbe03: y = 16'hfe00;
			16'hbe04: y = 16'hfe00;
			16'hbe05: y = 16'hfe00;
			16'hbe06: y = 16'hfe00;
			16'hbe07: y = 16'hfe00;
			16'hbe08: y = 16'hfe00;
			16'hbe09: y = 16'hfe00;
			16'hbe0a: y = 16'hfe00;
			16'hbe0b: y = 16'hfe00;
			16'hbe0c: y = 16'hfe00;
			16'hbe0d: y = 16'hfe00;
			16'hbe0e: y = 16'hfe00;
			16'hbe0f: y = 16'hfe00;
			16'hbe10: y = 16'hfe00;
			16'hbe11: y = 16'hfe00;
			16'hbe12: y = 16'hfe00;
			16'hbe13: y = 16'hfe00;
			16'hbe14: y = 16'hfe00;
			16'hbe15: y = 16'hfe00;
			16'hbe16: y = 16'hfe00;
			16'hbe17: y = 16'hfe00;
			16'hbe18: y = 16'hfe00;
			16'hbe19: y = 16'hfe00;
			16'hbe1a: y = 16'hfe00;
			16'hbe1b: y = 16'hfe00;
			16'hbe1c: y = 16'hfe00;
			16'hbe1d: y = 16'hfe00;
			16'hbe1e: y = 16'hfe00;
			16'hbe1f: y = 16'hfe00;
			16'hbe20: y = 16'hfe00;
			16'hbe21: y = 16'hfe00;
			16'hbe22: y = 16'hfe00;
			16'hbe23: y = 16'hfe00;
			16'hbe24: y = 16'hfe00;
			16'hbe25: y = 16'hfe00;
			16'hbe26: y = 16'hfe00;
			16'hbe27: y = 16'hfe00;
			16'hbe28: y = 16'hfe00;
			16'hbe29: y = 16'hfe00;
			16'hbe2a: y = 16'hfe00;
			16'hbe2b: y = 16'hfe00;
			16'hbe2c: y = 16'hfe00;
			16'hbe2d: y = 16'hfe00;
			16'hbe2e: y = 16'hfe00;
			16'hbe2f: y = 16'hfe00;
			16'hbe30: y = 16'hfe00;
			16'hbe31: y = 16'hfe00;
			16'hbe32: y = 16'hfe00;
			16'hbe33: y = 16'hfe00;
			16'hbe34: y = 16'hfe00;
			16'hbe35: y = 16'hfe00;
			16'hbe36: y = 16'hfe00;
			16'hbe37: y = 16'hfe00;
			16'hbe38: y = 16'hfe00;
			16'hbe39: y = 16'hfe00;
			16'hbe3a: y = 16'hfe00;
			16'hbe3b: y = 16'hfe00;
			16'hbe3c: y = 16'hfe00;
			16'hbe3d: y = 16'hfe00;
			16'hbe3e: y = 16'hfe00;
			16'hbe3f: y = 16'hfe00;
			16'hbe40: y = 16'hfe00;
			16'hbe41: y = 16'hfe00;
			16'hbe42: y = 16'hfe00;
			16'hbe43: y = 16'hfe00;
			16'hbe44: y = 16'hfe00;
			16'hbe45: y = 16'hfe00;
			16'hbe46: y = 16'hfe00;
			16'hbe47: y = 16'hfe00;
			16'hbe48: y = 16'hfe00;
			16'hbe49: y = 16'hfe00;
			16'hbe4a: y = 16'hfe00;
			16'hbe4b: y = 16'hfe00;
			16'hbe4c: y = 16'hfe00;
			16'hbe4d: y = 16'hfe00;
			16'hbe4e: y = 16'hfe00;
			16'hbe4f: y = 16'hfe00;
			16'hbe50: y = 16'hfe00;
			16'hbe51: y = 16'hfe00;
			16'hbe52: y = 16'hfe00;
			16'hbe53: y = 16'hfe00;
			16'hbe54: y = 16'hfe00;
			16'hbe55: y = 16'hfe00;
			16'hbe56: y = 16'hfe00;
			16'hbe57: y = 16'hfe00;
			16'hbe58: y = 16'hfe00;
			16'hbe59: y = 16'hfe00;
			16'hbe5a: y = 16'hfe00;
			16'hbe5b: y = 16'hfe00;
			16'hbe5c: y = 16'hfe00;
			16'hbe5d: y = 16'hfe00;
			16'hbe5e: y = 16'hfe00;
			16'hbe5f: y = 16'hfe00;
			16'hbe60: y = 16'hfe00;
			16'hbe61: y = 16'hfe00;
			16'hbe62: y = 16'hfe00;
			16'hbe63: y = 16'hfe00;
			16'hbe64: y = 16'hfe00;
			16'hbe65: y = 16'hfe00;
			16'hbe66: y = 16'hfe00;
			16'hbe67: y = 16'hfe00;
			16'hbe68: y = 16'hfe00;
			16'hbe69: y = 16'hfe00;
			16'hbe6a: y = 16'hfe00;
			16'hbe6b: y = 16'hfe00;
			16'hbe6c: y = 16'hfe00;
			16'hbe6d: y = 16'hfe00;
			16'hbe6e: y = 16'hfe00;
			16'hbe6f: y = 16'hfe00;
			16'hbe70: y = 16'hfe00;
			16'hbe71: y = 16'hfe00;
			16'hbe72: y = 16'hfe00;
			16'hbe73: y = 16'hfe00;
			16'hbe74: y = 16'hfe00;
			16'hbe75: y = 16'hfe00;
			16'hbe76: y = 16'hfe00;
			16'hbe77: y = 16'hfe00;
			16'hbe78: y = 16'hfe00;
			16'hbe79: y = 16'hfe00;
			16'hbe7a: y = 16'hfe00;
			16'hbe7b: y = 16'hfe00;
			16'hbe7c: y = 16'hfe00;
			16'hbe7d: y = 16'hfe00;
			16'hbe7e: y = 16'hfe00;
			16'hbe7f: y = 16'hfe00;
			16'hbe80: y = 16'hfe00;
			16'hbe81: y = 16'hfe00;
			16'hbe82: y = 16'hfe00;
			16'hbe83: y = 16'hfe00;
			16'hbe84: y = 16'hfe00;
			16'hbe85: y = 16'hfe00;
			16'hbe86: y = 16'hfe00;
			16'hbe87: y = 16'hfe00;
			16'hbe88: y = 16'hfe00;
			16'hbe89: y = 16'hfe00;
			16'hbe8a: y = 16'hfe00;
			16'hbe8b: y = 16'hfe00;
			16'hbe8c: y = 16'hfe00;
			16'hbe8d: y = 16'hfe00;
			16'hbe8e: y = 16'hfe00;
			16'hbe8f: y = 16'hfe00;
			16'hbe90: y = 16'hfe00;
			16'hbe91: y = 16'hfe00;
			16'hbe92: y = 16'hfe00;
			16'hbe93: y = 16'hfe00;
			16'hbe94: y = 16'hfe00;
			16'hbe95: y = 16'hfe00;
			16'hbe96: y = 16'hfe00;
			16'hbe97: y = 16'hfe00;
			16'hbe98: y = 16'hfe00;
			16'hbe99: y = 16'hfe00;
			16'hbe9a: y = 16'hfe00;
			16'hbe9b: y = 16'hfe00;
			16'hbe9c: y = 16'hfe00;
			16'hbe9d: y = 16'hfe00;
			16'hbe9e: y = 16'hfe00;
			16'hbe9f: y = 16'hfe00;
			16'hbea0: y = 16'hfe00;
			16'hbea1: y = 16'hfe00;
			16'hbea2: y = 16'hfe00;
			16'hbea3: y = 16'hfe00;
			16'hbea4: y = 16'hfe00;
			16'hbea5: y = 16'hfe00;
			16'hbea6: y = 16'hfe00;
			16'hbea7: y = 16'hfe00;
			16'hbea8: y = 16'hfe00;
			16'hbea9: y = 16'hfe00;
			16'hbeaa: y = 16'hfe00;
			16'hbeab: y = 16'hfe00;
			16'hbeac: y = 16'hfe00;
			16'hbead: y = 16'hfe00;
			16'hbeae: y = 16'hfe00;
			16'hbeaf: y = 16'hfe00;
			16'hbeb0: y = 16'hfe00;
			16'hbeb1: y = 16'hfe00;
			16'hbeb2: y = 16'hfe00;
			16'hbeb3: y = 16'hfe00;
			16'hbeb4: y = 16'hfe00;
			16'hbeb5: y = 16'hfe00;
			16'hbeb6: y = 16'hfe00;
			16'hbeb7: y = 16'hfe00;
			16'hbeb8: y = 16'hfe00;
			16'hbeb9: y = 16'hfe00;
			16'hbeba: y = 16'hfe00;
			16'hbebb: y = 16'hfe00;
			16'hbebc: y = 16'hfe00;
			16'hbebd: y = 16'hfe00;
			16'hbebe: y = 16'hfe00;
			16'hbebf: y = 16'hfe00;
			16'hbec0: y = 16'hfe00;
			16'hbec1: y = 16'hfe00;
			16'hbec2: y = 16'hfe00;
			16'hbec3: y = 16'hfe00;
			16'hbec4: y = 16'hfe00;
			16'hbec5: y = 16'hfe00;
			16'hbec6: y = 16'hfe00;
			16'hbec7: y = 16'hfe00;
			16'hbec8: y = 16'hfe00;
			16'hbec9: y = 16'hfe00;
			16'hbeca: y = 16'hfe00;
			16'hbecb: y = 16'hfe00;
			16'hbecc: y = 16'hfe00;
			16'hbecd: y = 16'hfe00;
			16'hbece: y = 16'hfe00;
			16'hbecf: y = 16'hfe00;
			16'hbed0: y = 16'hfe00;
			16'hbed1: y = 16'hfe00;
			16'hbed2: y = 16'hfe00;
			16'hbed3: y = 16'hfe00;
			16'hbed4: y = 16'hfe00;
			16'hbed5: y = 16'hfe00;
			16'hbed6: y = 16'hfe00;
			16'hbed7: y = 16'hfe00;
			16'hbed8: y = 16'hfe00;
			16'hbed9: y = 16'hfe00;
			16'hbeda: y = 16'hfe00;
			16'hbedb: y = 16'hfe00;
			16'hbedc: y = 16'hfe00;
			16'hbedd: y = 16'hfe00;
			16'hbede: y = 16'hfe00;
			16'hbedf: y = 16'hfe00;
			16'hbee0: y = 16'hfe00;
			16'hbee1: y = 16'hfe00;
			16'hbee2: y = 16'hfe00;
			16'hbee3: y = 16'hfe00;
			16'hbee4: y = 16'hfe00;
			16'hbee5: y = 16'hfe00;
			16'hbee6: y = 16'hfe00;
			16'hbee7: y = 16'hfe00;
			16'hbee8: y = 16'hfe00;
			16'hbee9: y = 16'hfe00;
			16'hbeea: y = 16'hfe00;
			16'hbeeb: y = 16'hfe00;
			16'hbeec: y = 16'hfe00;
			16'hbeed: y = 16'hfe00;
			16'hbeee: y = 16'hfe00;
			16'hbeef: y = 16'hfe00;
			16'hbef0: y = 16'hfe00;
			16'hbef1: y = 16'hfe00;
			16'hbef2: y = 16'hfe00;
			16'hbef3: y = 16'hfe00;
			16'hbef4: y = 16'hfe00;
			16'hbef5: y = 16'hfe00;
			16'hbef6: y = 16'hfe00;
			16'hbef7: y = 16'hfe00;
			16'hbef8: y = 16'hfe00;
			16'hbef9: y = 16'hfe00;
			16'hbefa: y = 16'hfe00;
			16'hbefb: y = 16'hfe00;
			16'hbefc: y = 16'hfe00;
			16'hbefd: y = 16'hfe00;
			16'hbefe: y = 16'hfe00;
			16'hbeff: y = 16'hfe00;
			16'hbf00: y = 16'hfe00;
			16'hbf01: y = 16'hfe00;
			16'hbf02: y = 16'hfe00;
			16'hbf03: y = 16'hfe00;
			16'hbf04: y = 16'hfe00;
			16'hbf05: y = 16'hfe00;
			16'hbf06: y = 16'hfe00;
			16'hbf07: y = 16'hfe00;
			16'hbf08: y = 16'hfe00;
			16'hbf09: y = 16'hfe00;
			16'hbf0a: y = 16'hfe00;
			16'hbf0b: y = 16'hfe00;
			16'hbf0c: y = 16'hfe00;
			16'hbf0d: y = 16'hfe00;
			16'hbf0e: y = 16'hfe00;
			16'hbf0f: y = 16'hfe00;
			16'hbf10: y = 16'hfe00;
			16'hbf11: y = 16'hfe00;
			16'hbf12: y = 16'hfe00;
			16'hbf13: y = 16'hfe00;
			16'hbf14: y = 16'hfe00;
			16'hbf15: y = 16'hfe00;
			16'hbf16: y = 16'hfe00;
			16'hbf17: y = 16'hfe00;
			16'hbf18: y = 16'hfe00;
			16'hbf19: y = 16'hfe00;
			16'hbf1a: y = 16'hfe00;
			16'hbf1b: y = 16'hfe00;
			16'hbf1c: y = 16'hfe00;
			16'hbf1d: y = 16'hfe00;
			16'hbf1e: y = 16'hfe00;
			16'hbf1f: y = 16'hfe00;
			16'hbf20: y = 16'hfe00;
			16'hbf21: y = 16'hfe00;
			16'hbf22: y = 16'hfe00;
			16'hbf23: y = 16'hfe00;
			16'hbf24: y = 16'hfe00;
			16'hbf25: y = 16'hfe00;
			16'hbf26: y = 16'hfe00;
			16'hbf27: y = 16'hfe00;
			16'hbf28: y = 16'hfe00;
			16'hbf29: y = 16'hfe00;
			16'hbf2a: y = 16'hfe00;
			16'hbf2b: y = 16'hfe00;
			16'hbf2c: y = 16'hfe00;
			16'hbf2d: y = 16'hfe00;
			16'hbf2e: y = 16'hfe00;
			16'hbf2f: y = 16'hfe00;
			16'hbf30: y = 16'hfe00;
			16'hbf31: y = 16'hfe00;
			16'hbf32: y = 16'hfe00;
			16'hbf33: y = 16'hfe00;
			16'hbf34: y = 16'hfe00;
			16'hbf35: y = 16'hfe00;
			16'hbf36: y = 16'hfe00;
			16'hbf37: y = 16'hfe00;
			16'hbf38: y = 16'hfe00;
			16'hbf39: y = 16'hfe00;
			16'hbf3a: y = 16'hfe00;
			16'hbf3b: y = 16'hfe00;
			16'hbf3c: y = 16'hfe00;
			16'hbf3d: y = 16'hfe00;
			16'hbf3e: y = 16'hfe00;
			16'hbf3f: y = 16'hfe00;
			16'hbf40: y = 16'hfe00;
			16'hbf41: y = 16'hfe00;
			16'hbf42: y = 16'hfe00;
			16'hbf43: y = 16'hfe00;
			16'hbf44: y = 16'hfe00;
			16'hbf45: y = 16'hfe00;
			16'hbf46: y = 16'hfe00;
			16'hbf47: y = 16'hfe00;
			16'hbf48: y = 16'hfe00;
			16'hbf49: y = 16'hfe00;
			16'hbf4a: y = 16'hfe00;
			16'hbf4b: y = 16'hfe00;
			16'hbf4c: y = 16'hfe00;
			16'hbf4d: y = 16'hfe00;
			16'hbf4e: y = 16'hfe00;
			16'hbf4f: y = 16'hfe00;
			16'hbf50: y = 16'hfe00;
			16'hbf51: y = 16'hfe00;
			16'hbf52: y = 16'hfe00;
			16'hbf53: y = 16'hfe00;
			16'hbf54: y = 16'hfe00;
			16'hbf55: y = 16'hfe00;
			16'hbf56: y = 16'hfe00;
			16'hbf57: y = 16'hfe00;
			16'hbf58: y = 16'hfe00;
			16'hbf59: y = 16'hfe00;
			16'hbf5a: y = 16'hfe00;
			16'hbf5b: y = 16'hfe00;
			16'hbf5c: y = 16'hfe00;
			16'hbf5d: y = 16'hfe00;
			16'hbf5e: y = 16'hfe00;
			16'hbf5f: y = 16'hfe00;
			16'hbf60: y = 16'hfe00;
			16'hbf61: y = 16'hfe00;
			16'hbf62: y = 16'hfe00;
			16'hbf63: y = 16'hfe00;
			16'hbf64: y = 16'hfe00;
			16'hbf65: y = 16'hfe00;
			16'hbf66: y = 16'hfe00;
			16'hbf67: y = 16'hfe00;
			16'hbf68: y = 16'hfe00;
			16'hbf69: y = 16'hfe00;
			16'hbf6a: y = 16'hfe00;
			16'hbf6b: y = 16'hfe00;
			16'hbf6c: y = 16'hfe00;
			16'hbf6d: y = 16'hfe00;
			16'hbf6e: y = 16'hfe00;
			16'hbf6f: y = 16'hfe00;
			16'hbf70: y = 16'hfe00;
			16'hbf71: y = 16'hfe00;
			16'hbf72: y = 16'hfe00;
			16'hbf73: y = 16'hfe00;
			16'hbf74: y = 16'hfe00;
			16'hbf75: y = 16'hfe00;
			16'hbf76: y = 16'hfe00;
			16'hbf77: y = 16'hfe00;
			16'hbf78: y = 16'hfe00;
			16'hbf79: y = 16'hfe00;
			16'hbf7a: y = 16'hfe00;
			16'hbf7b: y = 16'hfe00;
			16'hbf7c: y = 16'hfe00;
			16'hbf7d: y = 16'hfe00;
			16'hbf7e: y = 16'hfe00;
			16'hbf7f: y = 16'hfe00;
			16'hbf80: y = 16'hfe00;
			16'hbf81: y = 16'hfe00;
			16'hbf82: y = 16'hfe00;
			16'hbf83: y = 16'hfe00;
			16'hbf84: y = 16'hfe00;
			16'hbf85: y = 16'hfe00;
			16'hbf86: y = 16'hfe00;
			16'hbf87: y = 16'hfe00;
			16'hbf88: y = 16'hfe00;
			16'hbf89: y = 16'hfe00;
			16'hbf8a: y = 16'hfe00;
			16'hbf8b: y = 16'hfe00;
			16'hbf8c: y = 16'hfe00;
			16'hbf8d: y = 16'hfe00;
			16'hbf8e: y = 16'hfe00;
			16'hbf8f: y = 16'hfe00;
			16'hbf90: y = 16'hfe00;
			16'hbf91: y = 16'hfe00;
			16'hbf92: y = 16'hfe00;
			16'hbf93: y = 16'hfe00;
			16'hbf94: y = 16'hfe00;
			16'hbf95: y = 16'hfe00;
			16'hbf96: y = 16'hfe00;
			16'hbf97: y = 16'hfe00;
			16'hbf98: y = 16'hfe00;
			16'hbf99: y = 16'hfe00;
			16'hbf9a: y = 16'hfe00;
			16'hbf9b: y = 16'hfe00;
			16'hbf9c: y = 16'hfe00;
			16'hbf9d: y = 16'hfe00;
			16'hbf9e: y = 16'hfe00;
			16'hbf9f: y = 16'hfe00;
			16'hbfa0: y = 16'hfe00;
			16'hbfa1: y = 16'hfe00;
			16'hbfa2: y = 16'hfe00;
			16'hbfa3: y = 16'hfe00;
			16'hbfa4: y = 16'hfe00;
			16'hbfa5: y = 16'hfe00;
			16'hbfa6: y = 16'hfe00;
			16'hbfa7: y = 16'hfe00;
			16'hbfa8: y = 16'hfe00;
			16'hbfa9: y = 16'hfe00;
			16'hbfaa: y = 16'hfe00;
			16'hbfab: y = 16'hfe00;
			16'hbfac: y = 16'hfe00;
			16'hbfad: y = 16'hfe00;
			16'hbfae: y = 16'hfe00;
			16'hbfaf: y = 16'hfe00;
			16'hbfb0: y = 16'hfe00;
			16'hbfb1: y = 16'hfe00;
			16'hbfb2: y = 16'hfe00;
			16'hbfb3: y = 16'hfe00;
			16'hbfb4: y = 16'hfe00;
			16'hbfb5: y = 16'hfe00;
			16'hbfb6: y = 16'hfe00;
			16'hbfb7: y = 16'hfe00;
			16'hbfb8: y = 16'hfe00;
			16'hbfb9: y = 16'hfe00;
			16'hbfba: y = 16'hfe00;
			16'hbfbb: y = 16'hfe00;
			16'hbfbc: y = 16'hfe00;
			16'hbfbd: y = 16'hfe00;
			16'hbfbe: y = 16'hfe00;
			16'hbfbf: y = 16'hfe00;
			16'hbfc0: y = 16'hfe00;
			16'hbfc1: y = 16'hfe00;
			16'hbfc2: y = 16'hfe00;
			16'hbfc3: y = 16'hfe00;
			16'hbfc4: y = 16'hfe00;
			16'hbfc5: y = 16'hfe00;
			16'hbfc6: y = 16'hfe00;
			16'hbfc7: y = 16'hfe00;
			16'hbfc8: y = 16'hfe00;
			16'hbfc9: y = 16'hfe00;
			16'hbfca: y = 16'hfe00;
			16'hbfcb: y = 16'hfe00;
			16'hbfcc: y = 16'hfe00;
			16'hbfcd: y = 16'hfe00;
			16'hbfce: y = 16'hfe00;
			16'hbfcf: y = 16'hfe00;
			16'hbfd0: y = 16'hfe00;
			16'hbfd1: y = 16'hfe00;
			16'hbfd2: y = 16'hfe00;
			16'hbfd3: y = 16'hfe00;
			16'hbfd4: y = 16'hfe00;
			16'hbfd5: y = 16'hfe00;
			16'hbfd6: y = 16'hfe00;
			16'hbfd7: y = 16'hfe00;
			16'hbfd8: y = 16'hfe00;
			16'hbfd9: y = 16'hfe00;
			16'hbfda: y = 16'hfe00;
			16'hbfdb: y = 16'hfe00;
			16'hbfdc: y = 16'hfe00;
			16'hbfdd: y = 16'hfe00;
			16'hbfde: y = 16'hfe00;
			16'hbfdf: y = 16'hfe00;
			16'hbfe0: y = 16'hfe00;
			16'hbfe1: y = 16'hfe00;
			16'hbfe2: y = 16'hfe00;
			16'hbfe3: y = 16'hfe00;
			16'hbfe4: y = 16'hfe00;
			16'hbfe5: y = 16'hfe00;
			16'hbfe6: y = 16'hfe00;
			16'hbfe7: y = 16'hfe00;
			16'hbfe8: y = 16'hfe00;
			16'hbfe9: y = 16'hfe00;
			16'hbfea: y = 16'hfe00;
			16'hbfeb: y = 16'hfe00;
			16'hbfec: y = 16'hfe00;
			16'hbfed: y = 16'hfe00;
			16'hbfee: y = 16'hfe00;
			16'hbfef: y = 16'hfe00;
			16'hbff0: y = 16'hfe00;
			16'hbff1: y = 16'hfe00;
			16'hbff2: y = 16'hfe00;
			16'hbff3: y = 16'hfe00;
			16'hbff4: y = 16'hfe00;
			16'hbff5: y = 16'hfe00;
			16'hbff6: y = 16'hfe00;
			16'hbff7: y = 16'hfe00;
			16'hbff8: y = 16'hfe00;
			16'hbff9: y = 16'hfe00;
			16'hbffa: y = 16'hfe00;
			16'hbffb: y = 16'hfe00;
			16'hbffc: y = 16'hfe00;
			16'hbffd: y = 16'hfe00;
			16'hbffe: y = 16'hfe00;
			16'hbfff: y = 16'hfe00;
			16'hc000: y = 16'hfe00;
			16'hc001: y = 16'hfe00;
			16'hc002: y = 16'hfe00;
			16'hc003: y = 16'hfe00;
			16'hc004: y = 16'hfe00;
			16'hc005: y = 16'hfe00;
			16'hc006: y = 16'hfe00;
			16'hc007: y = 16'hfe00;
			16'hc008: y = 16'hfe00;
			16'hc009: y = 16'hfe00;
			16'hc00a: y = 16'hfe00;
			16'hc00b: y = 16'hfe00;
			16'hc00c: y = 16'hfe00;
			16'hc00d: y = 16'hfe00;
			16'hc00e: y = 16'hfe00;
			16'hc00f: y = 16'hfe00;
			16'hc010: y = 16'hfe00;
			16'hc011: y = 16'hfe00;
			16'hc012: y = 16'hfe00;
			16'hc013: y = 16'hfe00;
			16'hc014: y = 16'hfe00;
			16'hc015: y = 16'hfe00;
			16'hc016: y = 16'hfe00;
			16'hc017: y = 16'hfe00;
			16'hc018: y = 16'hfe00;
			16'hc019: y = 16'hfe00;
			16'hc01a: y = 16'hfe00;
			16'hc01b: y = 16'hfe00;
			16'hc01c: y = 16'hfe00;
			16'hc01d: y = 16'hfe00;
			16'hc01e: y = 16'hfe00;
			16'hc01f: y = 16'hfe00;
			16'hc020: y = 16'hfe00;
			16'hc021: y = 16'hfe00;
			16'hc022: y = 16'hfe00;
			16'hc023: y = 16'hfe00;
			16'hc024: y = 16'hfe00;
			16'hc025: y = 16'hfe00;
			16'hc026: y = 16'hfe00;
			16'hc027: y = 16'hfe00;
			16'hc028: y = 16'hfe00;
			16'hc029: y = 16'hfe00;
			16'hc02a: y = 16'hfe00;
			16'hc02b: y = 16'hfe00;
			16'hc02c: y = 16'hfe00;
			16'hc02d: y = 16'hfe00;
			16'hc02e: y = 16'hfe00;
			16'hc02f: y = 16'hfe00;
			16'hc030: y = 16'hfe00;
			16'hc031: y = 16'hfe00;
			16'hc032: y = 16'hfe00;
			16'hc033: y = 16'hfe00;
			16'hc034: y = 16'hfe00;
			16'hc035: y = 16'hfe00;
			16'hc036: y = 16'hfe00;
			16'hc037: y = 16'hfe00;
			16'hc038: y = 16'hfe00;
			16'hc039: y = 16'hfe00;
			16'hc03a: y = 16'hfe00;
			16'hc03b: y = 16'hfe00;
			16'hc03c: y = 16'hfe00;
			16'hc03d: y = 16'hfe00;
			16'hc03e: y = 16'hfe00;
			16'hc03f: y = 16'hfe00;
			16'hc040: y = 16'hfe00;
			16'hc041: y = 16'hfe00;
			16'hc042: y = 16'hfe00;
			16'hc043: y = 16'hfe00;
			16'hc044: y = 16'hfe00;
			16'hc045: y = 16'hfe00;
			16'hc046: y = 16'hfe00;
			16'hc047: y = 16'hfe00;
			16'hc048: y = 16'hfe00;
			16'hc049: y = 16'hfe00;
			16'hc04a: y = 16'hfe00;
			16'hc04b: y = 16'hfe00;
			16'hc04c: y = 16'hfe00;
			16'hc04d: y = 16'hfe00;
			16'hc04e: y = 16'hfe00;
			16'hc04f: y = 16'hfe00;
			16'hc050: y = 16'hfe00;
			16'hc051: y = 16'hfe00;
			16'hc052: y = 16'hfe00;
			16'hc053: y = 16'hfe00;
			16'hc054: y = 16'hfe00;
			16'hc055: y = 16'hfe00;
			16'hc056: y = 16'hfe00;
			16'hc057: y = 16'hfe00;
			16'hc058: y = 16'hfe00;
			16'hc059: y = 16'hfe00;
			16'hc05a: y = 16'hfe00;
			16'hc05b: y = 16'hfe00;
			16'hc05c: y = 16'hfe00;
			16'hc05d: y = 16'hfe00;
			16'hc05e: y = 16'hfe00;
			16'hc05f: y = 16'hfe00;
			16'hc060: y = 16'hfe00;
			16'hc061: y = 16'hfe00;
			16'hc062: y = 16'hfe00;
			16'hc063: y = 16'hfe00;
			16'hc064: y = 16'hfe00;
			16'hc065: y = 16'hfe00;
			16'hc066: y = 16'hfe00;
			16'hc067: y = 16'hfe00;
			16'hc068: y = 16'hfe00;
			16'hc069: y = 16'hfe00;
			16'hc06a: y = 16'hfe00;
			16'hc06b: y = 16'hfe00;
			16'hc06c: y = 16'hfe00;
			16'hc06d: y = 16'hfe00;
			16'hc06e: y = 16'hfe00;
			16'hc06f: y = 16'hfe00;
			16'hc070: y = 16'hfe00;
			16'hc071: y = 16'hfe00;
			16'hc072: y = 16'hfe00;
			16'hc073: y = 16'hfe00;
			16'hc074: y = 16'hfe00;
			16'hc075: y = 16'hfe00;
			16'hc076: y = 16'hfe00;
			16'hc077: y = 16'hfe00;
			16'hc078: y = 16'hfe00;
			16'hc079: y = 16'hfe00;
			16'hc07a: y = 16'hfe00;
			16'hc07b: y = 16'hfe00;
			16'hc07c: y = 16'hfe00;
			16'hc07d: y = 16'hfe00;
			16'hc07e: y = 16'hfe00;
			16'hc07f: y = 16'hfe00;
			16'hc080: y = 16'hfe00;
			16'hc081: y = 16'hfe00;
			16'hc082: y = 16'hfe00;
			16'hc083: y = 16'hfe00;
			16'hc084: y = 16'hfe00;
			16'hc085: y = 16'hfe00;
			16'hc086: y = 16'hfe00;
			16'hc087: y = 16'hfe00;
			16'hc088: y = 16'hfe00;
			16'hc089: y = 16'hfe00;
			16'hc08a: y = 16'hfe00;
			16'hc08b: y = 16'hfe00;
			16'hc08c: y = 16'hfe00;
			16'hc08d: y = 16'hfe00;
			16'hc08e: y = 16'hfe00;
			16'hc08f: y = 16'hfe00;
			16'hc090: y = 16'hfe00;
			16'hc091: y = 16'hfe00;
			16'hc092: y = 16'hfe00;
			16'hc093: y = 16'hfe00;
			16'hc094: y = 16'hfe00;
			16'hc095: y = 16'hfe00;
			16'hc096: y = 16'hfe00;
			16'hc097: y = 16'hfe00;
			16'hc098: y = 16'hfe00;
			16'hc099: y = 16'hfe00;
			16'hc09a: y = 16'hfe00;
			16'hc09b: y = 16'hfe00;
			16'hc09c: y = 16'hfe00;
			16'hc09d: y = 16'hfe00;
			16'hc09e: y = 16'hfe00;
			16'hc09f: y = 16'hfe00;
			16'hc0a0: y = 16'hfe00;
			16'hc0a1: y = 16'hfe00;
			16'hc0a2: y = 16'hfe00;
			16'hc0a3: y = 16'hfe00;
			16'hc0a4: y = 16'hfe00;
			16'hc0a5: y = 16'hfe00;
			16'hc0a6: y = 16'hfe00;
			16'hc0a7: y = 16'hfe00;
			16'hc0a8: y = 16'hfe00;
			16'hc0a9: y = 16'hfe00;
			16'hc0aa: y = 16'hfe00;
			16'hc0ab: y = 16'hfe00;
			16'hc0ac: y = 16'hfe00;
			16'hc0ad: y = 16'hfe00;
			16'hc0ae: y = 16'hfe00;
			16'hc0af: y = 16'hfe00;
			16'hc0b0: y = 16'hfe00;
			16'hc0b1: y = 16'hfe00;
			16'hc0b2: y = 16'hfe00;
			16'hc0b3: y = 16'hfe00;
			16'hc0b4: y = 16'hfe00;
			16'hc0b5: y = 16'hfe00;
			16'hc0b6: y = 16'hfe00;
			16'hc0b7: y = 16'hfe00;
			16'hc0b8: y = 16'hfe00;
			16'hc0b9: y = 16'hfe00;
			16'hc0ba: y = 16'hfe00;
			16'hc0bb: y = 16'hfe00;
			16'hc0bc: y = 16'hfe00;
			16'hc0bd: y = 16'hfe00;
			16'hc0be: y = 16'hfe00;
			16'hc0bf: y = 16'hfe00;
			16'hc0c0: y = 16'hfe00;
			16'hc0c1: y = 16'hfe00;
			16'hc0c2: y = 16'hfe00;
			16'hc0c3: y = 16'hfe00;
			16'hc0c4: y = 16'hfe00;
			16'hc0c5: y = 16'hfe00;
			16'hc0c6: y = 16'hfe00;
			16'hc0c7: y = 16'hfe00;
			16'hc0c8: y = 16'hfe00;
			16'hc0c9: y = 16'hfe00;
			16'hc0ca: y = 16'hfe00;
			16'hc0cb: y = 16'hfe00;
			16'hc0cc: y = 16'hfe00;
			16'hc0cd: y = 16'hfe00;
			16'hc0ce: y = 16'hfe00;
			16'hc0cf: y = 16'hfe00;
			16'hc0d0: y = 16'hfe00;
			16'hc0d1: y = 16'hfe00;
			16'hc0d2: y = 16'hfe00;
			16'hc0d3: y = 16'hfe00;
			16'hc0d4: y = 16'hfe00;
			16'hc0d5: y = 16'hfe00;
			16'hc0d6: y = 16'hfe00;
			16'hc0d7: y = 16'hfe00;
			16'hc0d8: y = 16'hfe00;
			16'hc0d9: y = 16'hfe00;
			16'hc0da: y = 16'hfe00;
			16'hc0db: y = 16'hfe00;
			16'hc0dc: y = 16'hfe00;
			16'hc0dd: y = 16'hfe00;
			16'hc0de: y = 16'hfe00;
			16'hc0df: y = 16'hfe00;
			16'hc0e0: y = 16'hfe00;
			16'hc0e1: y = 16'hfe00;
			16'hc0e2: y = 16'hfe00;
			16'hc0e3: y = 16'hfe00;
			16'hc0e4: y = 16'hfe00;
			16'hc0e5: y = 16'hfe00;
			16'hc0e6: y = 16'hfe00;
			16'hc0e7: y = 16'hfe00;
			16'hc0e8: y = 16'hfe00;
			16'hc0e9: y = 16'hfe00;
			16'hc0ea: y = 16'hfe00;
			16'hc0eb: y = 16'hfe00;
			16'hc0ec: y = 16'hfe00;
			16'hc0ed: y = 16'hfe00;
			16'hc0ee: y = 16'hfe00;
			16'hc0ef: y = 16'hfe00;
			16'hc0f0: y = 16'hfe00;
			16'hc0f1: y = 16'hfe00;
			16'hc0f2: y = 16'hfe00;
			16'hc0f3: y = 16'hfe00;
			16'hc0f4: y = 16'hfe00;
			16'hc0f5: y = 16'hfe00;
			16'hc0f6: y = 16'hfe00;
			16'hc0f7: y = 16'hfe00;
			16'hc0f8: y = 16'hfe00;
			16'hc0f9: y = 16'hfe00;
			16'hc0fa: y = 16'hfe00;
			16'hc0fb: y = 16'hfe00;
			16'hc0fc: y = 16'hfe00;
			16'hc0fd: y = 16'hfe00;
			16'hc0fe: y = 16'hfe00;
			16'hc0ff: y = 16'hfe00;
			16'hc100: y = 16'hfe00;
			16'hc101: y = 16'hfe00;
			16'hc102: y = 16'hfe00;
			16'hc103: y = 16'hfe00;
			16'hc104: y = 16'hfe00;
			16'hc105: y = 16'hfe00;
			16'hc106: y = 16'hfe00;
			16'hc107: y = 16'hfe00;
			16'hc108: y = 16'hfe00;
			16'hc109: y = 16'hfe00;
			16'hc10a: y = 16'hfe00;
			16'hc10b: y = 16'hfe00;
			16'hc10c: y = 16'hfe00;
			16'hc10d: y = 16'hfe00;
			16'hc10e: y = 16'hfe00;
			16'hc10f: y = 16'hfe00;
			16'hc110: y = 16'hfe00;
			16'hc111: y = 16'hfe00;
			16'hc112: y = 16'hfe00;
			16'hc113: y = 16'hfe00;
			16'hc114: y = 16'hfe00;
			16'hc115: y = 16'hfe00;
			16'hc116: y = 16'hfe00;
			16'hc117: y = 16'hfe00;
			16'hc118: y = 16'hfe00;
			16'hc119: y = 16'hfe00;
			16'hc11a: y = 16'hfe00;
			16'hc11b: y = 16'hfe00;
			16'hc11c: y = 16'hfe00;
			16'hc11d: y = 16'hfe00;
			16'hc11e: y = 16'hfe00;
			16'hc11f: y = 16'hfe00;
			16'hc120: y = 16'hfe00;
			16'hc121: y = 16'hfe00;
			16'hc122: y = 16'hfe00;
			16'hc123: y = 16'hfe00;
			16'hc124: y = 16'hfe00;
			16'hc125: y = 16'hfe00;
			16'hc126: y = 16'hfe00;
			16'hc127: y = 16'hfe00;
			16'hc128: y = 16'hfe00;
			16'hc129: y = 16'hfe00;
			16'hc12a: y = 16'hfe00;
			16'hc12b: y = 16'hfe00;
			16'hc12c: y = 16'hfe00;
			16'hc12d: y = 16'hfe00;
			16'hc12e: y = 16'hfe00;
			16'hc12f: y = 16'hfe00;
			16'hc130: y = 16'hfe00;
			16'hc131: y = 16'hfe00;
			16'hc132: y = 16'hfe00;
			16'hc133: y = 16'hfe00;
			16'hc134: y = 16'hfe00;
			16'hc135: y = 16'hfe00;
			16'hc136: y = 16'hfe00;
			16'hc137: y = 16'hfe00;
			16'hc138: y = 16'hfe00;
			16'hc139: y = 16'hfe00;
			16'hc13a: y = 16'hfe00;
			16'hc13b: y = 16'hfe00;
			16'hc13c: y = 16'hfe00;
			16'hc13d: y = 16'hfe00;
			16'hc13e: y = 16'hfe00;
			16'hc13f: y = 16'hfe00;
			16'hc140: y = 16'hfe00;
			16'hc141: y = 16'hfe00;
			16'hc142: y = 16'hfe00;
			16'hc143: y = 16'hfe00;
			16'hc144: y = 16'hfe00;
			16'hc145: y = 16'hfe00;
			16'hc146: y = 16'hfe00;
			16'hc147: y = 16'hfe00;
			16'hc148: y = 16'hfe00;
			16'hc149: y = 16'hfe00;
			16'hc14a: y = 16'hfe00;
			16'hc14b: y = 16'hfe00;
			16'hc14c: y = 16'hfe00;
			16'hc14d: y = 16'hfe00;
			16'hc14e: y = 16'hfe00;
			16'hc14f: y = 16'hfe00;
			16'hc150: y = 16'hfe00;
			16'hc151: y = 16'hfe00;
			16'hc152: y = 16'hfe00;
			16'hc153: y = 16'hfe00;
			16'hc154: y = 16'hfe00;
			16'hc155: y = 16'hfe00;
			16'hc156: y = 16'hfe00;
			16'hc157: y = 16'hfe00;
			16'hc158: y = 16'hfe00;
			16'hc159: y = 16'hfe00;
			16'hc15a: y = 16'hfe00;
			16'hc15b: y = 16'hfe00;
			16'hc15c: y = 16'hfe00;
			16'hc15d: y = 16'hfe00;
			16'hc15e: y = 16'hfe00;
			16'hc15f: y = 16'hfe00;
			16'hc160: y = 16'hfe00;
			16'hc161: y = 16'hfe00;
			16'hc162: y = 16'hfe00;
			16'hc163: y = 16'hfe00;
			16'hc164: y = 16'hfe00;
			16'hc165: y = 16'hfe00;
			16'hc166: y = 16'hfe00;
			16'hc167: y = 16'hfe00;
			16'hc168: y = 16'hfe00;
			16'hc169: y = 16'hfe00;
			16'hc16a: y = 16'hfe00;
			16'hc16b: y = 16'hfe00;
			16'hc16c: y = 16'hfe00;
			16'hc16d: y = 16'hfe00;
			16'hc16e: y = 16'hfe00;
			16'hc16f: y = 16'hfe00;
			16'hc170: y = 16'hfe00;
			16'hc171: y = 16'hfe00;
			16'hc172: y = 16'hfe00;
			16'hc173: y = 16'hfe00;
			16'hc174: y = 16'hfe00;
			16'hc175: y = 16'hfe00;
			16'hc176: y = 16'hfe00;
			16'hc177: y = 16'hfe00;
			16'hc178: y = 16'hfe00;
			16'hc179: y = 16'hfe00;
			16'hc17a: y = 16'hfe00;
			16'hc17b: y = 16'hfe00;
			16'hc17c: y = 16'hfe00;
			16'hc17d: y = 16'hfe00;
			16'hc17e: y = 16'hfe00;
			16'hc17f: y = 16'hfe00;
			16'hc180: y = 16'hfe00;
			16'hc181: y = 16'hfe00;
			16'hc182: y = 16'hfe00;
			16'hc183: y = 16'hfe00;
			16'hc184: y = 16'hfe00;
			16'hc185: y = 16'hfe00;
			16'hc186: y = 16'hfe00;
			16'hc187: y = 16'hfe00;
			16'hc188: y = 16'hfe00;
			16'hc189: y = 16'hfe00;
			16'hc18a: y = 16'hfe00;
			16'hc18b: y = 16'hfe00;
			16'hc18c: y = 16'hfe00;
			16'hc18d: y = 16'hfe00;
			16'hc18e: y = 16'hfe00;
			16'hc18f: y = 16'hfe00;
			16'hc190: y = 16'hfe00;
			16'hc191: y = 16'hfe00;
			16'hc192: y = 16'hfe00;
			16'hc193: y = 16'hfe00;
			16'hc194: y = 16'hfe00;
			16'hc195: y = 16'hfe00;
			16'hc196: y = 16'hfe00;
			16'hc197: y = 16'hfe00;
			16'hc198: y = 16'hfe00;
			16'hc199: y = 16'hfe00;
			16'hc19a: y = 16'hfe00;
			16'hc19b: y = 16'hfe00;
			16'hc19c: y = 16'hfe00;
			16'hc19d: y = 16'hfe00;
			16'hc19e: y = 16'hfe00;
			16'hc19f: y = 16'hfe00;
			16'hc1a0: y = 16'hfe00;
			16'hc1a1: y = 16'hfe00;
			16'hc1a2: y = 16'hfe00;
			16'hc1a3: y = 16'hfe00;
			16'hc1a4: y = 16'hfe00;
			16'hc1a5: y = 16'hfe00;
			16'hc1a6: y = 16'hfe00;
			16'hc1a7: y = 16'hfe00;
			16'hc1a8: y = 16'hfe00;
			16'hc1a9: y = 16'hfe00;
			16'hc1aa: y = 16'hfe00;
			16'hc1ab: y = 16'hfe00;
			16'hc1ac: y = 16'hfe00;
			16'hc1ad: y = 16'hfe00;
			16'hc1ae: y = 16'hfe00;
			16'hc1af: y = 16'hfe00;
			16'hc1b0: y = 16'hfe00;
			16'hc1b1: y = 16'hfe00;
			16'hc1b2: y = 16'hfe00;
			16'hc1b3: y = 16'hfe00;
			16'hc1b4: y = 16'hfe00;
			16'hc1b5: y = 16'hfe00;
			16'hc1b6: y = 16'hfe00;
			16'hc1b7: y = 16'hfe00;
			16'hc1b8: y = 16'hfe00;
			16'hc1b9: y = 16'hfe00;
			16'hc1ba: y = 16'hfe00;
			16'hc1bb: y = 16'hfe00;
			16'hc1bc: y = 16'hfe00;
			16'hc1bd: y = 16'hfe00;
			16'hc1be: y = 16'hfe00;
			16'hc1bf: y = 16'hfe00;
			16'hc1c0: y = 16'hfe00;
			16'hc1c1: y = 16'hfe00;
			16'hc1c2: y = 16'hfe00;
			16'hc1c3: y = 16'hfe00;
			16'hc1c4: y = 16'hfe00;
			16'hc1c5: y = 16'hfe00;
			16'hc1c6: y = 16'hfe00;
			16'hc1c7: y = 16'hfe00;
			16'hc1c8: y = 16'hfe00;
			16'hc1c9: y = 16'hfe00;
			16'hc1ca: y = 16'hfe00;
			16'hc1cb: y = 16'hfe00;
			16'hc1cc: y = 16'hfe00;
			16'hc1cd: y = 16'hfe00;
			16'hc1ce: y = 16'hfe00;
			16'hc1cf: y = 16'hfe00;
			16'hc1d0: y = 16'hfe00;
			16'hc1d1: y = 16'hfe00;
			16'hc1d2: y = 16'hfe00;
			16'hc1d3: y = 16'hfe00;
			16'hc1d4: y = 16'hfe00;
			16'hc1d5: y = 16'hfe00;
			16'hc1d6: y = 16'hfe00;
			16'hc1d7: y = 16'hfe00;
			16'hc1d8: y = 16'hfe00;
			16'hc1d9: y = 16'hfe00;
			16'hc1da: y = 16'hfe00;
			16'hc1db: y = 16'hfe00;
			16'hc1dc: y = 16'hfe00;
			16'hc1dd: y = 16'hfe00;
			16'hc1de: y = 16'hfe00;
			16'hc1df: y = 16'hfe00;
			16'hc1e0: y = 16'hfe00;
			16'hc1e1: y = 16'hfe00;
			16'hc1e2: y = 16'hfe00;
			16'hc1e3: y = 16'hfe00;
			16'hc1e4: y = 16'hfe00;
			16'hc1e5: y = 16'hfe00;
			16'hc1e6: y = 16'hfe00;
			16'hc1e7: y = 16'hfe00;
			16'hc1e8: y = 16'hfe00;
			16'hc1e9: y = 16'hfe00;
			16'hc1ea: y = 16'hfe00;
			16'hc1eb: y = 16'hfe00;
			16'hc1ec: y = 16'hfe00;
			16'hc1ed: y = 16'hfe00;
			16'hc1ee: y = 16'hfe00;
			16'hc1ef: y = 16'hfe00;
			16'hc1f0: y = 16'hfe00;
			16'hc1f1: y = 16'hfe00;
			16'hc1f2: y = 16'hfe00;
			16'hc1f3: y = 16'hfe00;
			16'hc1f4: y = 16'hfe00;
			16'hc1f5: y = 16'hfe00;
			16'hc1f6: y = 16'hfe00;
			16'hc1f7: y = 16'hfe00;
			16'hc1f8: y = 16'hfe00;
			16'hc1f9: y = 16'hfe00;
			16'hc1fa: y = 16'hfe00;
			16'hc1fb: y = 16'hfe00;
			16'hc1fc: y = 16'hfe00;
			16'hc1fd: y = 16'hfe00;
			16'hc1fe: y = 16'hfe00;
			16'hc1ff: y = 16'hfe00;
			16'hc200: y = 16'hfe00;
			16'hc201: y = 16'hfe00;
			16'hc202: y = 16'hfe00;
			16'hc203: y = 16'hfe00;
			16'hc204: y = 16'hfe00;
			16'hc205: y = 16'hfe00;
			16'hc206: y = 16'hfe00;
			16'hc207: y = 16'hfe00;
			16'hc208: y = 16'hfe00;
			16'hc209: y = 16'hfe00;
			16'hc20a: y = 16'hfe00;
			16'hc20b: y = 16'hfe00;
			16'hc20c: y = 16'hfe00;
			16'hc20d: y = 16'hfe00;
			16'hc20e: y = 16'hfe00;
			16'hc20f: y = 16'hfe00;
			16'hc210: y = 16'hfe00;
			16'hc211: y = 16'hfe00;
			16'hc212: y = 16'hfe00;
			16'hc213: y = 16'hfe00;
			16'hc214: y = 16'hfe00;
			16'hc215: y = 16'hfe00;
			16'hc216: y = 16'hfe00;
			16'hc217: y = 16'hfe00;
			16'hc218: y = 16'hfe00;
			16'hc219: y = 16'hfe00;
			16'hc21a: y = 16'hfe00;
			16'hc21b: y = 16'hfe00;
			16'hc21c: y = 16'hfe00;
			16'hc21d: y = 16'hfe00;
			16'hc21e: y = 16'hfe00;
			16'hc21f: y = 16'hfe00;
			16'hc220: y = 16'hfe00;
			16'hc221: y = 16'hfe00;
			16'hc222: y = 16'hfe00;
			16'hc223: y = 16'hfe00;
			16'hc224: y = 16'hfe00;
			16'hc225: y = 16'hfe00;
			16'hc226: y = 16'hfe00;
			16'hc227: y = 16'hfe00;
			16'hc228: y = 16'hfe00;
			16'hc229: y = 16'hfe00;
			16'hc22a: y = 16'hfe00;
			16'hc22b: y = 16'hfe00;
			16'hc22c: y = 16'hfe00;
			16'hc22d: y = 16'hfe00;
			16'hc22e: y = 16'hfe00;
			16'hc22f: y = 16'hfe00;
			16'hc230: y = 16'hfe00;
			16'hc231: y = 16'hfe00;
			16'hc232: y = 16'hfe00;
			16'hc233: y = 16'hfe00;
			16'hc234: y = 16'hfe00;
			16'hc235: y = 16'hfe00;
			16'hc236: y = 16'hfe00;
			16'hc237: y = 16'hfe00;
			16'hc238: y = 16'hfe00;
			16'hc239: y = 16'hfe00;
			16'hc23a: y = 16'hfe00;
			16'hc23b: y = 16'hfe00;
			16'hc23c: y = 16'hfe00;
			16'hc23d: y = 16'hfe00;
			16'hc23e: y = 16'hfe00;
			16'hc23f: y = 16'hfe00;
			16'hc240: y = 16'hfe00;
			16'hc241: y = 16'hfe00;
			16'hc242: y = 16'hfe00;
			16'hc243: y = 16'hfe00;
			16'hc244: y = 16'hfe00;
			16'hc245: y = 16'hfe00;
			16'hc246: y = 16'hfe00;
			16'hc247: y = 16'hfe00;
			16'hc248: y = 16'hfe00;
			16'hc249: y = 16'hfe00;
			16'hc24a: y = 16'hfe00;
			16'hc24b: y = 16'hfe00;
			16'hc24c: y = 16'hfe00;
			16'hc24d: y = 16'hfe00;
			16'hc24e: y = 16'hfe00;
			16'hc24f: y = 16'hfe00;
			16'hc250: y = 16'hfe00;
			16'hc251: y = 16'hfe00;
			16'hc252: y = 16'hfe00;
			16'hc253: y = 16'hfe00;
			16'hc254: y = 16'hfe00;
			16'hc255: y = 16'hfe00;
			16'hc256: y = 16'hfe00;
			16'hc257: y = 16'hfe00;
			16'hc258: y = 16'hfe00;
			16'hc259: y = 16'hfe00;
			16'hc25a: y = 16'hfe00;
			16'hc25b: y = 16'hfe00;
			16'hc25c: y = 16'hfe00;
			16'hc25d: y = 16'hfe00;
			16'hc25e: y = 16'hfe00;
			16'hc25f: y = 16'hfe00;
			16'hc260: y = 16'hfe00;
			16'hc261: y = 16'hfe00;
			16'hc262: y = 16'hfe00;
			16'hc263: y = 16'hfe00;
			16'hc264: y = 16'hfe00;
			16'hc265: y = 16'hfe00;
			16'hc266: y = 16'hfe00;
			16'hc267: y = 16'hfe00;
			16'hc268: y = 16'hfe00;
			16'hc269: y = 16'hfe00;
			16'hc26a: y = 16'hfe00;
			16'hc26b: y = 16'hfe00;
			16'hc26c: y = 16'hfe00;
			16'hc26d: y = 16'hfe00;
			16'hc26e: y = 16'hfe00;
			16'hc26f: y = 16'hfe00;
			16'hc270: y = 16'hfe00;
			16'hc271: y = 16'hfe00;
			16'hc272: y = 16'hfe00;
			16'hc273: y = 16'hfe00;
			16'hc274: y = 16'hfe00;
			16'hc275: y = 16'hfe00;
			16'hc276: y = 16'hfe00;
			16'hc277: y = 16'hfe00;
			16'hc278: y = 16'hfe00;
			16'hc279: y = 16'hfe00;
			16'hc27a: y = 16'hfe00;
			16'hc27b: y = 16'hfe00;
			16'hc27c: y = 16'hfe00;
			16'hc27d: y = 16'hfe00;
			16'hc27e: y = 16'hfe00;
			16'hc27f: y = 16'hfe00;
			16'hc280: y = 16'hfe00;
			16'hc281: y = 16'hfe00;
			16'hc282: y = 16'hfe00;
			16'hc283: y = 16'hfe00;
			16'hc284: y = 16'hfe00;
			16'hc285: y = 16'hfe00;
			16'hc286: y = 16'hfe00;
			16'hc287: y = 16'hfe00;
			16'hc288: y = 16'hfe00;
			16'hc289: y = 16'hfe00;
			16'hc28a: y = 16'hfe00;
			16'hc28b: y = 16'hfe00;
			16'hc28c: y = 16'hfe00;
			16'hc28d: y = 16'hfe00;
			16'hc28e: y = 16'hfe00;
			16'hc28f: y = 16'hfe00;
			16'hc290: y = 16'hfe00;
			16'hc291: y = 16'hfe00;
			16'hc292: y = 16'hfe00;
			16'hc293: y = 16'hfe00;
			16'hc294: y = 16'hfe00;
			16'hc295: y = 16'hfe00;
			16'hc296: y = 16'hfe00;
			16'hc297: y = 16'hfe00;
			16'hc298: y = 16'hfe00;
			16'hc299: y = 16'hfe00;
			16'hc29a: y = 16'hfe00;
			16'hc29b: y = 16'hfe00;
			16'hc29c: y = 16'hfe00;
			16'hc29d: y = 16'hfe00;
			16'hc29e: y = 16'hfe00;
			16'hc29f: y = 16'hfe00;
			16'hc2a0: y = 16'hfe00;
			16'hc2a1: y = 16'hfe00;
			16'hc2a2: y = 16'hfe00;
			16'hc2a3: y = 16'hfe00;
			16'hc2a4: y = 16'hfe00;
			16'hc2a5: y = 16'hfe00;
			16'hc2a6: y = 16'hfe00;
			16'hc2a7: y = 16'hfe00;
			16'hc2a8: y = 16'hfe00;
			16'hc2a9: y = 16'hfe00;
			16'hc2aa: y = 16'hfe00;
			16'hc2ab: y = 16'hfe00;
			16'hc2ac: y = 16'hfe00;
			16'hc2ad: y = 16'hfe00;
			16'hc2ae: y = 16'hfe00;
			16'hc2af: y = 16'hfe00;
			16'hc2b0: y = 16'hfe00;
			16'hc2b1: y = 16'hfe00;
			16'hc2b2: y = 16'hfe00;
			16'hc2b3: y = 16'hfe00;
			16'hc2b4: y = 16'hfe00;
			16'hc2b5: y = 16'hfe00;
			16'hc2b6: y = 16'hfe00;
			16'hc2b7: y = 16'hfe00;
			16'hc2b8: y = 16'hfe00;
			16'hc2b9: y = 16'hfe00;
			16'hc2ba: y = 16'hfe00;
			16'hc2bb: y = 16'hfe00;
			16'hc2bc: y = 16'hfe00;
			16'hc2bd: y = 16'hfe00;
			16'hc2be: y = 16'hfe00;
			16'hc2bf: y = 16'hfe00;
			16'hc2c0: y = 16'hfe00;
			16'hc2c1: y = 16'hfe00;
			16'hc2c2: y = 16'hfe00;
			16'hc2c3: y = 16'hfe00;
			16'hc2c4: y = 16'hfe00;
			16'hc2c5: y = 16'hfe00;
			16'hc2c6: y = 16'hfe00;
			16'hc2c7: y = 16'hfe00;
			16'hc2c8: y = 16'hfe00;
			16'hc2c9: y = 16'hfe00;
			16'hc2ca: y = 16'hfe00;
			16'hc2cb: y = 16'hfe00;
			16'hc2cc: y = 16'hfe00;
			16'hc2cd: y = 16'hfe00;
			16'hc2ce: y = 16'hfe00;
			16'hc2cf: y = 16'hfe00;
			16'hc2d0: y = 16'hfe00;
			16'hc2d1: y = 16'hfe00;
			16'hc2d2: y = 16'hfe00;
			16'hc2d3: y = 16'hfe00;
			16'hc2d4: y = 16'hfe00;
			16'hc2d5: y = 16'hfe00;
			16'hc2d6: y = 16'hfe00;
			16'hc2d7: y = 16'hfe00;
			16'hc2d8: y = 16'hfe00;
			16'hc2d9: y = 16'hfe00;
			16'hc2da: y = 16'hfe00;
			16'hc2db: y = 16'hfe00;
			16'hc2dc: y = 16'hfe00;
			16'hc2dd: y = 16'hfe00;
			16'hc2de: y = 16'hfe00;
			16'hc2df: y = 16'hfe00;
			16'hc2e0: y = 16'hfe00;
			16'hc2e1: y = 16'hfe00;
			16'hc2e2: y = 16'hfe00;
			16'hc2e3: y = 16'hfe00;
			16'hc2e4: y = 16'hfe00;
			16'hc2e5: y = 16'hfe00;
			16'hc2e6: y = 16'hfe00;
			16'hc2e7: y = 16'hfe00;
			16'hc2e8: y = 16'hfe00;
			16'hc2e9: y = 16'hfe00;
			16'hc2ea: y = 16'hfe00;
			16'hc2eb: y = 16'hfe00;
			16'hc2ec: y = 16'hfe00;
			16'hc2ed: y = 16'hfe00;
			16'hc2ee: y = 16'hfe00;
			16'hc2ef: y = 16'hfe00;
			16'hc2f0: y = 16'hfe00;
			16'hc2f1: y = 16'hfe00;
			16'hc2f2: y = 16'hfe00;
			16'hc2f3: y = 16'hfe00;
			16'hc2f4: y = 16'hfe00;
			16'hc2f5: y = 16'hfe00;
			16'hc2f6: y = 16'hfe00;
			16'hc2f7: y = 16'hfe00;
			16'hc2f8: y = 16'hfe00;
			16'hc2f9: y = 16'hfe00;
			16'hc2fa: y = 16'hfe00;
			16'hc2fb: y = 16'hfe00;
			16'hc2fc: y = 16'hfe00;
			16'hc2fd: y = 16'hfe00;
			16'hc2fe: y = 16'hfe00;
			16'hc2ff: y = 16'hfe00;
			16'hc300: y = 16'hfe00;
			16'hc301: y = 16'hfe00;
			16'hc302: y = 16'hfe00;
			16'hc303: y = 16'hfe00;
			16'hc304: y = 16'hfe00;
			16'hc305: y = 16'hfe00;
			16'hc306: y = 16'hfe00;
			16'hc307: y = 16'hfe00;
			16'hc308: y = 16'hfe00;
			16'hc309: y = 16'hfe00;
			16'hc30a: y = 16'hfe00;
			16'hc30b: y = 16'hfe00;
			16'hc30c: y = 16'hfe00;
			16'hc30d: y = 16'hfe00;
			16'hc30e: y = 16'hfe00;
			16'hc30f: y = 16'hfe00;
			16'hc310: y = 16'hfe00;
			16'hc311: y = 16'hfe00;
			16'hc312: y = 16'hfe00;
			16'hc313: y = 16'hfe00;
			16'hc314: y = 16'hfe00;
			16'hc315: y = 16'hfe00;
			16'hc316: y = 16'hfe00;
			16'hc317: y = 16'hfe00;
			16'hc318: y = 16'hfe00;
			16'hc319: y = 16'hfe00;
			16'hc31a: y = 16'hfe00;
			16'hc31b: y = 16'hfe00;
			16'hc31c: y = 16'hfe00;
			16'hc31d: y = 16'hfe00;
			16'hc31e: y = 16'hfe00;
			16'hc31f: y = 16'hfe00;
			16'hc320: y = 16'hfe00;
			16'hc321: y = 16'hfe00;
			16'hc322: y = 16'hfe00;
			16'hc323: y = 16'hfe00;
			16'hc324: y = 16'hfe00;
			16'hc325: y = 16'hfe00;
			16'hc326: y = 16'hfe00;
			16'hc327: y = 16'hfe00;
			16'hc328: y = 16'hfe00;
			16'hc329: y = 16'hfe00;
			16'hc32a: y = 16'hfe00;
			16'hc32b: y = 16'hfe00;
			16'hc32c: y = 16'hfe00;
			16'hc32d: y = 16'hfe00;
			16'hc32e: y = 16'hfe00;
			16'hc32f: y = 16'hfe00;
			16'hc330: y = 16'hfe00;
			16'hc331: y = 16'hfe00;
			16'hc332: y = 16'hfe00;
			16'hc333: y = 16'hfe00;
			16'hc334: y = 16'hfe00;
			16'hc335: y = 16'hfe00;
			16'hc336: y = 16'hfe00;
			16'hc337: y = 16'hfe00;
			16'hc338: y = 16'hfe00;
			16'hc339: y = 16'hfe00;
			16'hc33a: y = 16'hfe00;
			16'hc33b: y = 16'hfe00;
			16'hc33c: y = 16'hfe00;
			16'hc33d: y = 16'hfe00;
			16'hc33e: y = 16'hfe00;
			16'hc33f: y = 16'hfe00;
			16'hc340: y = 16'hfe00;
			16'hc341: y = 16'hfe00;
			16'hc342: y = 16'hfe00;
			16'hc343: y = 16'hfe00;
			16'hc344: y = 16'hfe00;
			16'hc345: y = 16'hfe00;
			16'hc346: y = 16'hfe00;
			16'hc347: y = 16'hfe00;
			16'hc348: y = 16'hfe00;
			16'hc349: y = 16'hfe00;
			16'hc34a: y = 16'hfe00;
			16'hc34b: y = 16'hfe00;
			16'hc34c: y = 16'hfe00;
			16'hc34d: y = 16'hfe00;
			16'hc34e: y = 16'hfe00;
			16'hc34f: y = 16'hfe00;
			16'hc350: y = 16'hfe00;
			16'hc351: y = 16'hfe00;
			16'hc352: y = 16'hfe00;
			16'hc353: y = 16'hfe00;
			16'hc354: y = 16'hfe00;
			16'hc355: y = 16'hfe00;
			16'hc356: y = 16'hfe00;
			16'hc357: y = 16'hfe00;
			16'hc358: y = 16'hfe00;
			16'hc359: y = 16'hfe00;
			16'hc35a: y = 16'hfe00;
			16'hc35b: y = 16'hfe00;
			16'hc35c: y = 16'hfe00;
			16'hc35d: y = 16'hfe00;
			16'hc35e: y = 16'hfe00;
			16'hc35f: y = 16'hfe00;
			16'hc360: y = 16'hfe00;
			16'hc361: y = 16'hfe00;
			16'hc362: y = 16'hfe00;
			16'hc363: y = 16'hfe00;
			16'hc364: y = 16'hfe00;
			16'hc365: y = 16'hfe00;
			16'hc366: y = 16'hfe00;
			16'hc367: y = 16'hfe00;
			16'hc368: y = 16'hfe00;
			16'hc369: y = 16'hfe00;
			16'hc36a: y = 16'hfe00;
			16'hc36b: y = 16'hfe00;
			16'hc36c: y = 16'hfe00;
			16'hc36d: y = 16'hfe00;
			16'hc36e: y = 16'hfe00;
			16'hc36f: y = 16'hfe00;
			16'hc370: y = 16'hfe00;
			16'hc371: y = 16'hfe00;
			16'hc372: y = 16'hfe00;
			16'hc373: y = 16'hfe00;
			16'hc374: y = 16'hfe00;
			16'hc375: y = 16'hfe00;
			16'hc376: y = 16'hfe00;
			16'hc377: y = 16'hfe00;
			16'hc378: y = 16'hfe00;
			16'hc379: y = 16'hfe00;
			16'hc37a: y = 16'hfe00;
			16'hc37b: y = 16'hfe00;
			16'hc37c: y = 16'hfe00;
			16'hc37d: y = 16'hfe00;
			16'hc37e: y = 16'hfe00;
			16'hc37f: y = 16'hfe00;
			16'hc380: y = 16'hfe00;
			16'hc381: y = 16'hfe00;
			16'hc382: y = 16'hfe00;
			16'hc383: y = 16'hfe00;
			16'hc384: y = 16'hfe00;
			16'hc385: y = 16'hfe00;
			16'hc386: y = 16'hfe00;
			16'hc387: y = 16'hfe00;
			16'hc388: y = 16'hfe00;
			16'hc389: y = 16'hfe00;
			16'hc38a: y = 16'hfe00;
			16'hc38b: y = 16'hfe00;
			16'hc38c: y = 16'hfe00;
			16'hc38d: y = 16'hfe00;
			16'hc38e: y = 16'hfe00;
			16'hc38f: y = 16'hfe00;
			16'hc390: y = 16'hfe00;
			16'hc391: y = 16'hfe00;
			16'hc392: y = 16'hfe00;
			16'hc393: y = 16'hfe00;
			16'hc394: y = 16'hfe00;
			16'hc395: y = 16'hfe00;
			16'hc396: y = 16'hfe00;
			16'hc397: y = 16'hfe00;
			16'hc398: y = 16'hfe00;
			16'hc399: y = 16'hfe00;
			16'hc39a: y = 16'hfe00;
			16'hc39b: y = 16'hfe00;
			16'hc39c: y = 16'hfe00;
			16'hc39d: y = 16'hfe00;
			16'hc39e: y = 16'hfe00;
			16'hc39f: y = 16'hfe00;
			16'hc3a0: y = 16'hfe00;
			16'hc3a1: y = 16'hfe00;
			16'hc3a2: y = 16'hfe00;
			16'hc3a3: y = 16'hfe00;
			16'hc3a4: y = 16'hfe00;
			16'hc3a5: y = 16'hfe00;
			16'hc3a6: y = 16'hfe00;
			16'hc3a7: y = 16'hfe00;
			16'hc3a8: y = 16'hfe00;
			16'hc3a9: y = 16'hfe00;
			16'hc3aa: y = 16'hfe00;
			16'hc3ab: y = 16'hfe00;
			16'hc3ac: y = 16'hfe00;
			16'hc3ad: y = 16'hfe00;
			16'hc3ae: y = 16'hfe00;
			16'hc3af: y = 16'hfe00;
			16'hc3b0: y = 16'hfe00;
			16'hc3b1: y = 16'hfe00;
			16'hc3b2: y = 16'hfe00;
			16'hc3b3: y = 16'hfe00;
			16'hc3b4: y = 16'hfe00;
			16'hc3b5: y = 16'hfe00;
			16'hc3b6: y = 16'hfe00;
			16'hc3b7: y = 16'hfe00;
			16'hc3b8: y = 16'hfe00;
			16'hc3b9: y = 16'hfe00;
			16'hc3ba: y = 16'hfe00;
			16'hc3bb: y = 16'hfe00;
			16'hc3bc: y = 16'hfe00;
			16'hc3bd: y = 16'hfe00;
			16'hc3be: y = 16'hfe00;
			16'hc3bf: y = 16'hfe00;
			16'hc3c0: y = 16'hfe00;
			16'hc3c1: y = 16'hfe00;
			16'hc3c2: y = 16'hfe00;
			16'hc3c3: y = 16'hfe00;
			16'hc3c4: y = 16'hfe00;
			16'hc3c5: y = 16'hfe00;
			16'hc3c6: y = 16'hfe00;
			16'hc3c7: y = 16'hfe00;
			16'hc3c8: y = 16'hfe00;
			16'hc3c9: y = 16'hfe00;
			16'hc3ca: y = 16'hfe00;
			16'hc3cb: y = 16'hfe00;
			16'hc3cc: y = 16'hfe00;
			16'hc3cd: y = 16'hfe00;
			16'hc3ce: y = 16'hfe00;
			16'hc3cf: y = 16'hfe00;
			16'hc3d0: y = 16'hfe00;
			16'hc3d1: y = 16'hfe00;
			16'hc3d2: y = 16'hfe00;
			16'hc3d3: y = 16'hfe00;
			16'hc3d4: y = 16'hfe00;
			16'hc3d5: y = 16'hfe00;
			16'hc3d6: y = 16'hfe00;
			16'hc3d7: y = 16'hfe00;
			16'hc3d8: y = 16'hfe00;
			16'hc3d9: y = 16'hfe00;
			16'hc3da: y = 16'hfe00;
			16'hc3db: y = 16'hfe00;
			16'hc3dc: y = 16'hfe00;
			16'hc3dd: y = 16'hfe00;
			16'hc3de: y = 16'hfe00;
			16'hc3df: y = 16'hfe00;
			16'hc3e0: y = 16'hfe00;
			16'hc3e1: y = 16'hfe00;
			16'hc3e2: y = 16'hfe00;
			16'hc3e3: y = 16'hfe00;
			16'hc3e4: y = 16'hfe00;
			16'hc3e5: y = 16'hfe00;
			16'hc3e6: y = 16'hfe00;
			16'hc3e7: y = 16'hfe00;
			16'hc3e8: y = 16'hfe00;
			16'hc3e9: y = 16'hfe00;
			16'hc3ea: y = 16'hfe00;
			16'hc3eb: y = 16'hfe00;
			16'hc3ec: y = 16'hfe00;
			16'hc3ed: y = 16'hfe00;
			16'hc3ee: y = 16'hfe00;
			16'hc3ef: y = 16'hfe00;
			16'hc3f0: y = 16'hfe00;
			16'hc3f1: y = 16'hfe00;
			16'hc3f2: y = 16'hfe00;
			16'hc3f3: y = 16'hfe00;
			16'hc3f4: y = 16'hfe00;
			16'hc3f5: y = 16'hfe00;
			16'hc3f6: y = 16'hfe00;
			16'hc3f7: y = 16'hfe00;
			16'hc3f8: y = 16'hfe00;
			16'hc3f9: y = 16'hfe00;
			16'hc3fa: y = 16'hfe00;
			16'hc3fb: y = 16'hfe00;
			16'hc3fc: y = 16'hfe00;
			16'hc3fd: y = 16'hfe00;
			16'hc3fe: y = 16'hfe00;
			16'hc3ff: y = 16'hfe00;
			16'hc400: y = 16'hfe00;
			16'hc401: y = 16'hfe00;
			16'hc402: y = 16'hfe00;
			16'hc403: y = 16'hfe00;
			16'hc404: y = 16'hfe00;
			16'hc405: y = 16'hfe00;
			16'hc406: y = 16'hfe00;
			16'hc407: y = 16'hfe00;
			16'hc408: y = 16'hfe00;
			16'hc409: y = 16'hfe00;
			16'hc40a: y = 16'hfe00;
			16'hc40b: y = 16'hfe00;
			16'hc40c: y = 16'hfe00;
			16'hc40d: y = 16'hfe00;
			16'hc40e: y = 16'hfe00;
			16'hc40f: y = 16'hfe00;
			16'hc410: y = 16'hfe00;
			16'hc411: y = 16'hfe00;
			16'hc412: y = 16'hfe00;
			16'hc413: y = 16'hfe00;
			16'hc414: y = 16'hfe00;
			16'hc415: y = 16'hfe00;
			16'hc416: y = 16'hfe00;
			16'hc417: y = 16'hfe00;
			16'hc418: y = 16'hfe00;
			16'hc419: y = 16'hfe00;
			16'hc41a: y = 16'hfe00;
			16'hc41b: y = 16'hfe00;
			16'hc41c: y = 16'hfe00;
			16'hc41d: y = 16'hfe00;
			16'hc41e: y = 16'hfe00;
			16'hc41f: y = 16'hfe00;
			16'hc420: y = 16'hfe00;
			16'hc421: y = 16'hfe00;
			16'hc422: y = 16'hfe00;
			16'hc423: y = 16'hfe00;
			16'hc424: y = 16'hfe00;
			16'hc425: y = 16'hfe00;
			16'hc426: y = 16'hfe00;
			16'hc427: y = 16'hfe00;
			16'hc428: y = 16'hfe00;
			16'hc429: y = 16'hfe00;
			16'hc42a: y = 16'hfe00;
			16'hc42b: y = 16'hfe00;
			16'hc42c: y = 16'hfe00;
			16'hc42d: y = 16'hfe00;
			16'hc42e: y = 16'hfe00;
			16'hc42f: y = 16'hfe00;
			16'hc430: y = 16'hfe00;
			16'hc431: y = 16'hfe00;
			16'hc432: y = 16'hfe00;
			16'hc433: y = 16'hfe00;
			16'hc434: y = 16'hfe00;
			16'hc435: y = 16'hfe00;
			16'hc436: y = 16'hfe00;
			16'hc437: y = 16'hfe00;
			16'hc438: y = 16'hfe00;
			16'hc439: y = 16'hfe00;
			16'hc43a: y = 16'hfe00;
			16'hc43b: y = 16'hfe00;
			16'hc43c: y = 16'hfe00;
			16'hc43d: y = 16'hfe00;
			16'hc43e: y = 16'hfe00;
			16'hc43f: y = 16'hfe00;
			16'hc440: y = 16'hfe00;
			16'hc441: y = 16'hfe00;
			16'hc442: y = 16'hfe00;
			16'hc443: y = 16'hfe00;
			16'hc444: y = 16'hfe00;
			16'hc445: y = 16'hfe00;
			16'hc446: y = 16'hfe00;
			16'hc447: y = 16'hfe00;
			16'hc448: y = 16'hfe00;
			16'hc449: y = 16'hfe00;
			16'hc44a: y = 16'hfe00;
			16'hc44b: y = 16'hfe00;
			16'hc44c: y = 16'hfe00;
			16'hc44d: y = 16'hfe00;
			16'hc44e: y = 16'hfe00;
			16'hc44f: y = 16'hfe00;
			16'hc450: y = 16'hfe00;
			16'hc451: y = 16'hfe00;
			16'hc452: y = 16'hfe00;
			16'hc453: y = 16'hfe00;
			16'hc454: y = 16'hfe00;
			16'hc455: y = 16'hfe00;
			16'hc456: y = 16'hfe00;
			16'hc457: y = 16'hfe00;
			16'hc458: y = 16'hfe00;
			16'hc459: y = 16'hfe00;
			16'hc45a: y = 16'hfe00;
			16'hc45b: y = 16'hfe00;
			16'hc45c: y = 16'hfe00;
			16'hc45d: y = 16'hfe00;
			16'hc45e: y = 16'hfe00;
			16'hc45f: y = 16'hfe00;
			16'hc460: y = 16'hfe00;
			16'hc461: y = 16'hfe00;
			16'hc462: y = 16'hfe00;
			16'hc463: y = 16'hfe00;
			16'hc464: y = 16'hfe00;
			16'hc465: y = 16'hfe00;
			16'hc466: y = 16'hfe00;
			16'hc467: y = 16'hfe00;
			16'hc468: y = 16'hfe00;
			16'hc469: y = 16'hfe00;
			16'hc46a: y = 16'hfe00;
			16'hc46b: y = 16'hfe00;
			16'hc46c: y = 16'hfe00;
			16'hc46d: y = 16'hfe00;
			16'hc46e: y = 16'hfe00;
			16'hc46f: y = 16'hfe00;
			16'hc470: y = 16'hfe00;
			16'hc471: y = 16'hfe00;
			16'hc472: y = 16'hfe00;
			16'hc473: y = 16'hfe00;
			16'hc474: y = 16'hfe00;
			16'hc475: y = 16'hfe00;
			16'hc476: y = 16'hfe00;
			16'hc477: y = 16'hfe00;
			16'hc478: y = 16'hfe00;
			16'hc479: y = 16'hfe00;
			16'hc47a: y = 16'hfe00;
			16'hc47b: y = 16'hfe00;
			16'hc47c: y = 16'hfe00;
			16'hc47d: y = 16'hfe00;
			16'hc47e: y = 16'hfe00;
			16'hc47f: y = 16'hfe00;
			16'hc480: y = 16'hfe00;
			16'hc481: y = 16'hfe00;
			16'hc482: y = 16'hfe00;
			16'hc483: y = 16'hfe00;
			16'hc484: y = 16'hfe00;
			16'hc485: y = 16'hfe00;
			16'hc486: y = 16'hfe00;
			16'hc487: y = 16'hfe00;
			16'hc488: y = 16'hfe00;
			16'hc489: y = 16'hfe00;
			16'hc48a: y = 16'hfe00;
			16'hc48b: y = 16'hfe00;
			16'hc48c: y = 16'hfe00;
			16'hc48d: y = 16'hfe00;
			16'hc48e: y = 16'hfe00;
			16'hc48f: y = 16'hfe00;
			16'hc490: y = 16'hfe00;
			16'hc491: y = 16'hfe00;
			16'hc492: y = 16'hfe00;
			16'hc493: y = 16'hfe00;
			16'hc494: y = 16'hfe00;
			16'hc495: y = 16'hfe00;
			16'hc496: y = 16'hfe00;
			16'hc497: y = 16'hfe00;
			16'hc498: y = 16'hfe00;
			16'hc499: y = 16'hfe00;
			16'hc49a: y = 16'hfe00;
			16'hc49b: y = 16'hfe00;
			16'hc49c: y = 16'hfe00;
			16'hc49d: y = 16'hfe00;
			16'hc49e: y = 16'hfe00;
			16'hc49f: y = 16'hfe00;
			16'hc4a0: y = 16'hfe00;
			16'hc4a1: y = 16'hfe00;
			16'hc4a2: y = 16'hfe00;
			16'hc4a3: y = 16'hfe00;
			16'hc4a4: y = 16'hfe00;
			16'hc4a5: y = 16'hfe00;
			16'hc4a6: y = 16'hfe00;
			16'hc4a7: y = 16'hfe00;
			16'hc4a8: y = 16'hfe00;
			16'hc4a9: y = 16'hfe00;
			16'hc4aa: y = 16'hfe00;
			16'hc4ab: y = 16'hfe00;
			16'hc4ac: y = 16'hfe00;
			16'hc4ad: y = 16'hfe00;
			16'hc4ae: y = 16'hfe00;
			16'hc4af: y = 16'hfe00;
			16'hc4b0: y = 16'hfe00;
			16'hc4b1: y = 16'hfe00;
			16'hc4b2: y = 16'hfe00;
			16'hc4b3: y = 16'hfe00;
			16'hc4b4: y = 16'hfe00;
			16'hc4b5: y = 16'hfe00;
			16'hc4b6: y = 16'hfe00;
			16'hc4b7: y = 16'hfe00;
			16'hc4b8: y = 16'hfe00;
			16'hc4b9: y = 16'hfe00;
			16'hc4ba: y = 16'hfe00;
			16'hc4bb: y = 16'hfe00;
			16'hc4bc: y = 16'hfe00;
			16'hc4bd: y = 16'hfe00;
			16'hc4be: y = 16'hfe00;
			16'hc4bf: y = 16'hfe00;
			16'hc4c0: y = 16'hfe00;
			16'hc4c1: y = 16'hfe00;
			16'hc4c2: y = 16'hfe00;
			16'hc4c3: y = 16'hfe00;
			16'hc4c4: y = 16'hfe00;
			16'hc4c5: y = 16'hfe00;
			16'hc4c6: y = 16'hfe00;
			16'hc4c7: y = 16'hfe00;
			16'hc4c8: y = 16'hfe00;
			16'hc4c9: y = 16'hfe00;
			16'hc4ca: y = 16'hfe00;
			16'hc4cb: y = 16'hfe00;
			16'hc4cc: y = 16'hfe00;
			16'hc4cd: y = 16'hfe00;
			16'hc4ce: y = 16'hfe00;
			16'hc4cf: y = 16'hfe00;
			16'hc4d0: y = 16'hfe00;
			16'hc4d1: y = 16'hfe00;
			16'hc4d2: y = 16'hfe00;
			16'hc4d3: y = 16'hfe00;
			16'hc4d4: y = 16'hfe00;
			16'hc4d5: y = 16'hfe00;
			16'hc4d6: y = 16'hfe00;
			16'hc4d7: y = 16'hfe00;
			16'hc4d8: y = 16'hfe00;
			16'hc4d9: y = 16'hfe00;
			16'hc4da: y = 16'hfe00;
			16'hc4db: y = 16'hfe00;
			16'hc4dc: y = 16'hfe00;
			16'hc4dd: y = 16'hfe00;
			16'hc4de: y = 16'hfe00;
			16'hc4df: y = 16'hfe00;
			16'hc4e0: y = 16'hfe00;
			16'hc4e1: y = 16'hfe00;
			16'hc4e2: y = 16'hfe00;
			16'hc4e3: y = 16'hfe00;
			16'hc4e4: y = 16'hfe00;
			16'hc4e5: y = 16'hfe00;
			16'hc4e6: y = 16'hfe00;
			16'hc4e7: y = 16'hfe00;
			16'hc4e8: y = 16'hfe00;
			16'hc4e9: y = 16'hfe00;
			16'hc4ea: y = 16'hfe00;
			16'hc4eb: y = 16'hfe00;
			16'hc4ec: y = 16'hfe00;
			16'hc4ed: y = 16'hfe00;
			16'hc4ee: y = 16'hfe00;
			16'hc4ef: y = 16'hfe00;
			16'hc4f0: y = 16'hfe00;
			16'hc4f1: y = 16'hfe00;
			16'hc4f2: y = 16'hfe00;
			16'hc4f3: y = 16'hfe00;
			16'hc4f4: y = 16'hfe00;
			16'hc4f5: y = 16'hfe00;
			16'hc4f6: y = 16'hfe00;
			16'hc4f7: y = 16'hfe00;
			16'hc4f8: y = 16'hfe00;
			16'hc4f9: y = 16'hfe00;
			16'hc4fa: y = 16'hfe00;
			16'hc4fb: y = 16'hfe00;
			16'hc4fc: y = 16'hfe00;
			16'hc4fd: y = 16'hfe00;
			16'hc4fe: y = 16'hfe00;
			16'hc4ff: y = 16'hfe00;
			16'hc500: y = 16'hfe00;
			16'hc501: y = 16'hfe00;
			16'hc502: y = 16'hfe00;
			16'hc503: y = 16'hfe00;
			16'hc504: y = 16'hfe00;
			16'hc505: y = 16'hfe00;
			16'hc506: y = 16'hfe00;
			16'hc507: y = 16'hfe00;
			16'hc508: y = 16'hfe00;
			16'hc509: y = 16'hfe00;
			16'hc50a: y = 16'hfe00;
			16'hc50b: y = 16'hfe00;
			16'hc50c: y = 16'hfe00;
			16'hc50d: y = 16'hfe00;
			16'hc50e: y = 16'hfe00;
			16'hc50f: y = 16'hfe00;
			16'hc510: y = 16'hfe00;
			16'hc511: y = 16'hfe00;
			16'hc512: y = 16'hfe00;
			16'hc513: y = 16'hfe00;
			16'hc514: y = 16'hfe00;
			16'hc515: y = 16'hfe00;
			16'hc516: y = 16'hfe00;
			16'hc517: y = 16'hfe00;
			16'hc518: y = 16'hfe00;
			16'hc519: y = 16'hfe00;
			16'hc51a: y = 16'hfe00;
			16'hc51b: y = 16'hfe00;
			16'hc51c: y = 16'hfe00;
			16'hc51d: y = 16'hfe00;
			16'hc51e: y = 16'hfe00;
			16'hc51f: y = 16'hfe00;
			16'hc520: y = 16'hfe00;
			16'hc521: y = 16'hfe00;
			16'hc522: y = 16'hfe00;
			16'hc523: y = 16'hfe00;
			16'hc524: y = 16'hfe00;
			16'hc525: y = 16'hfe00;
			16'hc526: y = 16'hfe00;
			16'hc527: y = 16'hfe00;
			16'hc528: y = 16'hfe00;
			16'hc529: y = 16'hfe00;
			16'hc52a: y = 16'hfe00;
			16'hc52b: y = 16'hfe00;
			16'hc52c: y = 16'hfe00;
			16'hc52d: y = 16'hfe00;
			16'hc52e: y = 16'hfe00;
			16'hc52f: y = 16'hfe00;
			16'hc530: y = 16'hfe00;
			16'hc531: y = 16'hfe00;
			16'hc532: y = 16'hfe00;
			16'hc533: y = 16'hfe00;
			16'hc534: y = 16'hfe00;
			16'hc535: y = 16'hfe00;
			16'hc536: y = 16'hfe00;
			16'hc537: y = 16'hfe00;
			16'hc538: y = 16'hfe00;
			16'hc539: y = 16'hfe00;
			16'hc53a: y = 16'hfe00;
			16'hc53b: y = 16'hfe00;
			16'hc53c: y = 16'hfe00;
			16'hc53d: y = 16'hfe00;
			16'hc53e: y = 16'hfe00;
			16'hc53f: y = 16'hfe00;
			16'hc540: y = 16'hfe00;
			16'hc541: y = 16'hfe00;
			16'hc542: y = 16'hfe00;
			16'hc543: y = 16'hfe00;
			16'hc544: y = 16'hfe00;
			16'hc545: y = 16'hfe00;
			16'hc546: y = 16'hfe00;
			16'hc547: y = 16'hfe00;
			16'hc548: y = 16'hfe00;
			16'hc549: y = 16'hfe00;
			16'hc54a: y = 16'hfe00;
			16'hc54b: y = 16'hfe00;
			16'hc54c: y = 16'hfe00;
			16'hc54d: y = 16'hfe00;
			16'hc54e: y = 16'hfe00;
			16'hc54f: y = 16'hfe00;
			16'hc550: y = 16'hfe00;
			16'hc551: y = 16'hfe00;
			16'hc552: y = 16'hfe00;
			16'hc553: y = 16'hfe00;
			16'hc554: y = 16'hfe00;
			16'hc555: y = 16'hfe00;
			16'hc556: y = 16'hfe00;
			16'hc557: y = 16'hfe00;
			16'hc558: y = 16'hfe00;
			16'hc559: y = 16'hfe00;
			16'hc55a: y = 16'hfe00;
			16'hc55b: y = 16'hfe00;
			16'hc55c: y = 16'hfe00;
			16'hc55d: y = 16'hfe00;
			16'hc55e: y = 16'hfe00;
			16'hc55f: y = 16'hfe00;
			16'hc560: y = 16'hfe00;
			16'hc561: y = 16'hfe00;
			16'hc562: y = 16'hfe00;
			16'hc563: y = 16'hfe00;
			16'hc564: y = 16'hfe00;
			16'hc565: y = 16'hfe00;
			16'hc566: y = 16'hfe00;
			16'hc567: y = 16'hfe00;
			16'hc568: y = 16'hfe00;
			16'hc569: y = 16'hfe00;
			16'hc56a: y = 16'hfe00;
			16'hc56b: y = 16'hfe00;
			16'hc56c: y = 16'hfe00;
			16'hc56d: y = 16'hfe00;
			16'hc56e: y = 16'hfe00;
			16'hc56f: y = 16'hfe00;
			16'hc570: y = 16'hfe00;
			16'hc571: y = 16'hfe00;
			16'hc572: y = 16'hfe00;
			16'hc573: y = 16'hfe00;
			16'hc574: y = 16'hfe00;
			16'hc575: y = 16'hfe00;
			16'hc576: y = 16'hfe00;
			16'hc577: y = 16'hfe00;
			16'hc578: y = 16'hfe00;
			16'hc579: y = 16'hfe00;
			16'hc57a: y = 16'hfe00;
			16'hc57b: y = 16'hfe00;
			16'hc57c: y = 16'hfe00;
			16'hc57d: y = 16'hfe00;
			16'hc57e: y = 16'hfe00;
			16'hc57f: y = 16'hfe00;
			16'hc580: y = 16'hfe00;
			16'hc581: y = 16'hfe00;
			16'hc582: y = 16'hfe00;
			16'hc583: y = 16'hfe00;
			16'hc584: y = 16'hfe00;
			16'hc585: y = 16'hfe00;
			16'hc586: y = 16'hfe00;
			16'hc587: y = 16'hfe00;
			16'hc588: y = 16'hfe00;
			16'hc589: y = 16'hfe00;
			16'hc58a: y = 16'hfe00;
			16'hc58b: y = 16'hfe00;
			16'hc58c: y = 16'hfe00;
			16'hc58d: y = 16'hfe00;
			16'hc58e: y = 16'hfe00;
			16'hc58f: y = 16'hfe00;
			16'hc590: y = 16'hfe00;
			16'hc591: y = 16'hfe00;
			16'hc592: y = 16'hfe00;
			16'hc593: y = 16'hfe00;
			16'hc594: y = 16'hfe00;
			16'hc595: y = 16'hfe00;
			16'hc596: y = 16'hfe00;
			16'hc597: y = 16'hfe00;
			16'hc598: y = 16'hfe00;
			16'hc599: y = 16'hfe00;
			16'hc59a: y = 16'hfe00;
			16'hc59b: y = 16'hfe00;
			16'hc59c: y = 16'hfe00;
			16'hc59d: y = 16'hfe00;
			16'hc59e: y = 16'hfe00;
			16'hc59f: y = 16'hfe00;
			16'hc5a0: y = 16'hfe00;
			16'hc5a1: y = 16'hfe00;
			16'hc5a2: y = 16'hfe00;
			16'hc5a3: y = 16'hfe00;
			16'hc5a4: y = 16'hfe00;
			16'hc5a5: y = 16'hfe00;
			16'hc5a6: y = 16'hfe00;
			16'hc5a7: y = 16'hfe00;
			16'hc5a8: y = 16'hfe00;
			16'hc5a9: y = 16'hfe00;
			16'hc5aa: y = 16'hfe00;
			16'hc5ab: y = 16'hfe00;
			16'hc5ac: y = 16'hfe00;
			16'hc5ad: y = 16'hfe00;
			16'hc5ae: y = 16'hfe00;
			16'hc5af: y = 16'hfe00;
			16'hc5b0: y = 16'hfe00;
			16'hc5b1: y = 16'hfe00;
			16'hc5b2: y = 16'hfe00;
			16'hc5b3: y = 16'hfe00;
			16'hc5b4: y = 16'hfe00;
			16'hc5b5: y = 16'hfe00;
			16'hc5b6: y = 16'hfe00;
			16'hc5b7: y = 16'hfe00;
			16'hc5b8: y = 16'hfe00;
			16'hc5b9: y = 16'hfe00;
			16'hc5ba: y = 16'hfe00;
			16'hc5bb: y = 16'hfe00;
			16'hc5bc: y = 16'hfe00;
			16'hc5bd: y = 16'hfe00;
			16'hc5be: y = 16'hfe00;
			16'hc5bf: y = 16'hfe00;
			16'hc5c0: y = 16'hfe00;
			16'hc5c1: y = 16'hfe00;
			16'hc5c2: y = 16'hfe00;
			16'hc5c3: y = 16'hfe00;
			16'hc5c4: y = 16'hfe00;
			16'hc5c5: y = 16'hfe00;
			16'hc5c6: y = 16'hfe00;
			16'hc5c7: y = 16'hfe00;
			16'hc5c8: y = 16'hfe00;
			16'hc5c9: y = 16'hfe00;
			16'hc5ca: y = 16'hfe00;
			16'hc5cb: y = 16'hfe00;
			16'hc5cc: y = 16'hfe00;
			16'hc5cd: y = 16'hfe00;
			16'hc5ce: y = 16'hfe00;
			16'hc5cf: y = 16'hfe00;
			16'hc5d0: y = 16'hfe00;
			16'hc5d1: y = 16'hfe00;
			16'hc5d2: y = 16'hfe00;
			16'hc5d3: y = 16'hfe00;
			16'hc5d4: y = 16'hfe00;
			16'hc5d5: y = 16'hfe00;
			16'hc5d6: y = 16'hfe00;
			16'hc5d7: y = 16'hfe00;
			16'hc5d8: y = 16'hfe00;
			16'hc5d9: y = 16'hfe00;
			16'hc5da: y = 16'hfe00;
			16'hc5db: y = 16'hfe00;
			16'hc5dc: y = 16'hfe00;
			16'hc5dd: y = 16'hfe00;
			16'hc5de: y = 16'hfe00;
			16'hc5df: y = 16'hfe00;
			16'hc5e0: y = 16'hfe00;
			16'hc5e1: y = 16'hfe00;
			16'hc5e2: y = 16'hfe00;
			16'hc5e3: y = 16'hfe00;
			16'hc5e4: y = 16'hfe00;
			16'hc5e5: y = 16'hfe00;
			16'hc5e6: y = 16'hfe00;
			16'hc5e7: y = 16'hfe00;
			16'hc5e8: y = 16'hfe00;
			16'hc5e9: y = 16'hfe00;
			16'hc5ea: y = 16'hfe00;
			16'hc5eb: y = 16'hfe00;
			16'hc5ec: y = 16'hfe00;
			16'hc5ed: y = 16'hfe00;
			16'hc5ee: y = 16'hfe00;
			16'hc5ef: y = 16'hfe00;
			16'hc5f0: y = 16'hfe00;
			16'hc5f1: y = 16'hfe00;
			16'hc5f2: y = 16'hfe00;
			16'hc5f3: y = 16'hfe00;
			16'hc5f4: y = 16'hfe00;
			16'hc5f5: y = 16'hfe00;
			16'hc5f6: y = 16'hfe00;
			16'hc5f7: y = 16'hfe00;
			16'hc5f8: y = 16'hfe00;
			16'hc5f9: y = 16'hfe00;
			16'hc5fa: y = 16'hfe00;
			16'hc5fb: y = 16'hfe00;
			16'hc5fc: y = 16'hfe00;
			16'hc5fd: y = 16'hfe00;
			16'hc5fe: y = 16'hfe00;
			16'hc5ff: y = 16'hfe00;
			16'hc600: y = 16'hfe00;
			16'hc601: y = 16'hfe00;
			16'hc602: y = 16'hfe00;
			16'hc603: y = 16'hfe00;
			16'hc604: y = 16'hfe00;
			16'hc605: y = 16'hfe00;
			16'hc606: y = 16'hfe00;
			16'hc607: y = 16'hfe00;
			16'hc608: y = 16'hfe00;
			16'hc609: y = 16'hfe00;
			16'hc60a: y = 16'hfe00;
			16'hc60b: y = 16'hfe00;
			16'hc60c: y = 16'hfe00;
			16'hc60d: y = 16'hfe00;
			16'hc60e: y = 16'hfe00;
			16'hc60f: y = 16'hfe00;
			16'hc610: y = 16'hfe00;
			16'hc611: y = 16'hfe00;
			16'hc612: y = 16'hfe00;
			16'hc613: y = 16'hfe00;
			16'hc614: y = 16'hfe00;
			16'hc615: y = 16'hfe00;
			16'hc616: y = 16'hfe00;
			16'hc617: y = 16'hfe00;
			16'hc618: y = 16'hfe00;
			16'hc619: y = 16'hfe00;
			16'hc61a: y = 16'hfe00;
			16'hc61b: y = 16'hfe00;
			16'hc61c: y = 16'hfe00;
			16'hc61d: y = 16'hfe00;
			16'hc61e: y = 16'hfe00;
			16'hc61f: y = 16'hfe00;
			16'hc620: y = 16'hfe00;
			16'hc621: y = 16'hfe00;
			16'hc622: y = 16'hfe00;
			16'hc623: y = 16'hfe00;
			16'hc624: y = 16'hfe00;
			16'hc625: y = 16'hfe00;
			16'hc626: y = 16'hfe00;
			16'hc627: y = 16'hfe00;
			16'hc628: y = 16'hfe00;
			16'hc629: y = 16'hfe00;
			16'hc62a: y = 16'hfe00;
			16'hc62b: y = 16'hfe00;
			16'hc62c: y = 16'hfe00;
			16'hc62d: y = 16'hfe00;
			16'hc62e: y = 16'hfe00;
			16'hc62f: y = 16'hfe00;
			16'hc630: y = 16'hfe00;
			16'hc631: y = 16'hfe00;
			16'hc632: y = 16'hfe00;
			16'hc633: y = 16'hfe00;
			16'hc634: y = 16'hfe00;
			16'hc635: y = 16'hfe00;
			16'hc636: y = 16'hfe00;
			16'hc637: y = 16'hfe00;
			16'hc638: y = 16'hfe00;
			16'hc639: y = 16'hfe00;
			16'hc63a: y = 16'hfe00;
			16'hc63b: y = 16'hfe00;
			16'hc63c: y = 16'hfe00;
			16'hc63d: y = 16'hfe00;
			16'hc63e: y = 16'hfe00;
			16'hc63f: y = 16'hfe00;
			16'hc640: y = 16'hfe00;
			16'hc641: y = 16'hfe00;
			16'hc642: y = 16'hfe00;
			16'hc643: y = 16'hfe00;
			16'hc644: y = 16'hfe00;
			16'hc645: y = 16'hfe00;
			16'hc646: y = 16'hfe00;
			16'hc647: y = 16'hfe00;
			16'hc648: y = 16'hfe00;
			16'hc649: y = 16'hfe00;
			16'hc64a: y = 16'hfe00;
			16'hc64b: y = 16'hfe00;
			16'hc64c: y = 16'hfe00;
			16'hc64d: y = 16'hfe00;
			16'hc64e: y = 16'hfe00;
			16'hc64f: y = 16'hfe00;
			16'hc650: y = 16'hfe00;
			16'hc651: y = 16'hfe00;
			16'hc652: y = 16'hfe00;
			16'hc653: y = 16'hfe00;
			16'hc654: y = 16'hfe00;
			16'hc655: y = 16'hfe00;
			16'hc656: y = 16'hfe00;
			16'hc657: y = 16'hfe00;
			16'hc658: y = 16'hfe00;
			16'hc659: y = 16'hfe00;
			16'hc65a: y = 16'hfe00;
			16'hc65b: y = 16'hfe00;
			16'hc65c: y = 16'hfe00;
			16'hc65d: y = 16'hfe00;
			16'hc65e: y = 16'hfe00;
			16'hc65f: y = 16'hfe00;
			16'hc660: y = 16'hfe00;
			16'hc661: y = 16'hfe00;
			16'hc662: y = 16'hfe00;
			16'hc663: y = 16'hfe00;
			16'hc664: y = 16'hfe00;
			16'hc665: y = 16'hfe00;
			16'hc666: y = 16'hfe00;
			16'hc667: y = 16'hfe00;
			16'hc668: y = 16'hfe00;
			16'hc669: y = 16'hfe00;
			16'hc66a: y = 16'hfe00;
			16'hc66b: y = 16'hfe00;
			16'hc66c: y = 16'hfe00;
			16'hc66d: y = 16'hfe00;
			16'hc66e: y = 16'hfe00;
			16'hc66f: y = 16'hfe00;
			16'hc670: y = 16'hfe00;
			16'hc671: y = 16'hfe00;
			16'hc672: y = 16'hfe00;
			16'hc673: y = 16'hfe00;
			16'hc674: y = 16'hfe00;
			16'hc675: y = 16'hfe00;
			16'hc676: y = 16'hfe00;
			16'hc677: y = 16'hfe00;
			16'hc678: y = 16'hfe00;
			16'hc679: y = 16'hfe00;
			16'hc67a: y = 16'hfe00;
			16'hc67b: y = 16'hfe00;
			16'hc67c: y = 16'hfe00;
			16'hc67d: y = 16'hfe00;
			16'hc67e: y = 16'hfe00;
			16'hc67f: y = 16'hfe00;
			16'hc680: y = 16'hfe00;
			16'hc681: y = 16'hfe00;
			16'hc682: y = 16'hfe00;
			16'hc683: y = 16'hfe00;
			16'hc684: y = 16'hfe00;
			16'hc685: y = 16'hfe00;
			16'hc686: y = 16'hfe00;
			16'hc687: y = 16'hfe00;
			16'hc688: y = 16'hfe00;
			16'hc689: y = 16'hfe00;
			16'hc68a: y = 16'hfe00;
			16'hc68b: y = 16'hfe00;
			16'hc68c: y = 16'hfe00;
			16'hc68d: y = 16'hfe00;
			16'hc68e: y = 16'hfe00;
			16'hc68f: y = 16'hfe00;
			16'hc690: y = 16'hfe00;
			16'hc691: y = 16'hfe00;
			16'hc692: y = 16'hfe00;
			16'hc693: y = 16'hfe00;
			16'hc694: y = 16'hfe00;
			16'hc695: y = 16'hfe00;
			16'hc696: y = 16'hfe00;
			16'hc697: y = 16'hfe00;
			16'hc698: y = 16'hfe00;
			16'hc699: y = 16'hfe00;
			16'hc69a: y = 16'hfe00;
			16'hc69b: y = 16'hfe00;
			16'hc69c: y = 16'hfe00;
			16'hc69d: y = 16'hfe00;
			16'hc69e: y = 16'hfe00;
			16'hc69f: y = 16'hfe00;
			16'hc6a0: y = 16'hfe00;
			16'hc6a1: y = 16'hfe00;
			16'hc6a2: y = 16'hfe00;
			16'hc6a3: y = 16'hfe00;
			16'hc6a4: y = 16'hfe00;
			16'hc6a5: y = 16'hfe00;
			16'hc6a6: y = 16'hfe00;
			16'hc6a7: y = 16'hfe00;
			16'hc6a8: y = 16'hfe00;
			16'hc6a9: y = 16'hfe00;
			16'hc6aa: y = 16'hfe00;
			16'hc6ab: y = 16'hfe00;
			16'hc6ac: y = 16'hfe00;
			16'hc6ad: y = 16'hfe00;
			16'hc6ae: y = 16'hfe00;
			16'hc6af: y = 16'hfe00;
			16'hc6b0: y = 16'hfe00;
			16'hc6b1: y = 16'hfe00;
			16'hc6b2: y = 16'hfe00;
			16'hc6b3: y = 16'hfe00;
			16'hc6b4: y = 16'hfe00;
			16'hc6b5: y = 16'hfe00;
			16'hc6b6: y = 16'hfe00;
			16'hc6b7: y = 16'hfe00;
			16'hc6b8: y = 16'hfe00;
			16'hc6b9: y = 16'hfe00;
			16'hc6ba: y = 16'hfe00;
			16'hc6bb: y = 16'hfe00;
			16'hc6bc: y = 16'hfe00;
			16'hc6bd: y = 16'hfe00;
			16'hc6be: y = 16'hfe00;
			16'hc6bf: y = 16'hfe00;
			16'hc6c0: y = 16'hfe00;
			16'hc6c1: y = 16'hfe00;
			16'hc6c2: y = 16'hfe00;
			16'hc6c3: y = 16'hfe00;
			16'hc6c4: y = 16'hfe00;
			16'hc6c5: y = 16'hfe00;
			16'hc6c6: y = 16'hfe00;
			16'hc6c7: y = 16'hfe00;
			16'hc6c8: y = 16'hfe00;
			16'hc6c9: y = 16'hfe00;
			16'hc6ca: y = 16'hfe00;
			16'hc6cb: y = 16'hfe00;
			16'hc6cc: y = 16'hfe00;
			16'hc6cd: y = 16'hfe00;
			16'hc6ce: y = 16'hfe00;
			16'hc6cf: y = 16'hfe00;
			16'hc6d0: y = 16'hfe00;
			16'hc6d1: y = 16'hfe00;
			16'hc6d2: y = 16'hfe00;
			16'hc6d3: y = 16'hfe00;
			16'hc6d4: y = 16'hfe00;
			16'hc6d5: y = 16'hfe00;
			16'hc6d6: y = 16'hfe00;
			16'hc6d7: y = 16'hfe00;
			16'hc6d8: y = 16'hfe00;
			16'hc6d9: y = 16'hfe00;
			16'hc6da: y = 16'hfe00;
			16'hc6db: y = 16'hfe00;
			16'hc6dc: y = 16'hfe00;
			16'hc6dd: y = 16'hfe00;
			16'hc6de: y = 16'hfe00;
			16'hc6df: y = 16'hfe00;
			16'hc6e0: y = 16'hfe00;
			16'hc6e1: y = 16'hfe00;
			16'hc6e2: y = 16'hfe00;
			16'hc6e3: y = 16'hfe00;
			16'hc6e4: y = 16'hfe00;
			16'hc6e5: y = 16'hfe00;
			16'hc6e6: y = 16'hfe00;
			16'hc6e7: y = 16'hfe00;
			16'hc6e8: y = 16'hfe00;
			16'hc6e9: y = 16'hfe00;
			16'hc6ea: y = 16'hfe00;
			16'hc6eb: y = 16'hfe00;
			16'hc6ec: y = 16'hfe00;
			16'hc6ed: y = 16'hfe00;
			16'hc6ee: y = 16'hfe00;
			16'hc6ef: y = 16'hfe00;
			16'hc6f0: y = 16'hfe00;
			16'hc6f1: y = 16'hfe00;
			16'hc6f2: y = 16'hfe00;
			16'hc6f3: y = 16'hfe00;
			16'hc6f4: y = 16'hfe00;
			16'hc6f5: y = 16'hfe00;
			16'hc6f6: y = 16'hfe00;
			16'hc6f7: y = 16'hfe00;
			16'hc6f8: y = 16'hfe00;
			16'hc6f9: y = 16'hfe00;
			16'hc6fa: y = 16'hfe00;
			16'hc6fb: y = 16'hfe00;
			16'hc6fc: y = 16'hfe00;
			16'hc6fd: y = 16'hfe00;
			16'hc6fe: y = 16'hfe00;
			16'hc6ff: y = 16'hfe00;
			16'hc700: y = 16'hfe00;
			16'hc701: y = 16'hfe00;
			16'hc702: y = 16'hfe00;
			16'hc703: y = 16'hfe00;
			16'hc704: y = 16'hfe00;
			16'hc705: y = 16'hfe00;
			16'hc706: y = 16'hfe00;
			16'hc707: y = 16'hfe00;
			16'hc708: y = 16'hfe00;
			16'hc709: y = 16'hfe00;
			16'hc70a: y = 16'hfe00;
			16'hc70b: y = 16'hfe00;
			16'hc70c: y = 16'hfe00;
			16'hc70d: y = 16'hfe00;
			16'hc70e: y = 16'hfe00;
			16'hc70f: y = 16'hfe00;
			16'hc710: y = 16'hfe00;
			16'hc711: y = 16'hfe00;
			16'hc712: y = 16'hfe00;
			16'hc713: y = 16'hfe00;
			16'hc714: y = 16'hfe00;
			16'hc715: y = 16'hfe00;
			16'hc716: y = 16'hfe00;
			16'hc717: y = 16'hfe00;
			16'hc718: y = 16'hfe00;
			16'hc719: y = 16'hfe00;
			16'hc71a: y = 16'hfe00;
			16'hc71b: y = 16'hfe00;
			16'hc71c: y = 16'hfe00;
			16'hc71d: y = 16'hfe00;
			16'hc71e: y = 16'hfe00;
			16'hc71f: y = 16'hfe00;
			16'hc720: y = 16'hfe00;
			16'hc721: y = 16'hfe00;
			16'hc722: y = 16'hfe00;
			16'hc723: y = 16'hfe00;
			16'hc724: y = 16'hfe00;
			16'hc725: y = 16'hfe00;
			16'hc726: y = 16'hfe00;
			16'hc727: y = 16'hfe00;
			16'hc728: y = 16'hfe00;
			16'hc729: y = 16'hfe00;
			16'hc72a: y = 16'hfe00;
			16'hc72b: y = 16'hfe00;
			16'hc72c: y = 16'hfe00;
			16'hc72d: y = 16'hfe00;
			16'hc72e: y = 16'hfe00;
			16'hc72f: y = 16'hfe00;
			16'hc730: y = 16'hfe00;
			16'hc731: y = 16'hfe00;
			16'hc732: y = 16'hfe00;
			16'hc733: y = 16'hfe00;
			16'hc734: y = 16'hfe00;
			16'hc735: y = 16'hfe00;
			16'hc736: y = 16'hfe00;
			16'hc737: y = 16'hfe00;
			16'hc738: y = 16'hfe00;
			16'hc739: y = 16'hfe00;
			16'hc73a: y = 16'hfe00;
			16'hc73b: y = 16'hfe00;
			16'hc73c: y = 16'hfe00;
			16'hc73d: y = 16'hfe00;
			16'hc73e: y = 16'hfe00;
			16'hc73f: y = 16'hfe00;
			16'hc740: y = 16'hfe00;
			16'hc741: y = 16'hfe00;
			16'hc742: y = 16'hfe00;
			16'hc743: y = 16'hfe00;
			16'hc744: y = 16'hfe00;
			16'hc745: y = 16'hfe00;
			16'hc746: y = 16'hfe00;
			16'hc747: y = 16'hfe00;
			16'hc748: y = 16'hfe00;
			16'hc749: y = 16'hfe00;
			16'hc74a: y = 16'hfe00;
			16'hc74b: y = 16'hfe00;
			16'hc74c: y = 16'hfe00;
			16'hc74d: y = 16'hfe00;
			16'hc74e: y = 16'hfe00;
			16'hc74f: y = 16'hfe00;
			16'hc750: y = 16'hfe00;
			16'hc751: y = 16'hfe00;
			16'hc752: y = 16'hfe00;
			16'hc753: y = 16'hfe00;
			16'hc754: y = 16'hfe00;
			16'hc755: y = 16'hfe00;
			16'hc756: y = 16'hfe00;
			16'hc757: y = 16'hfe00;
			16'hc758: y = 16'hfe00;
			16'hc759: y = 16'hfe00;
			16'hc75a: y = 16'hfe00;
			16'hc75b: y = 16'hfe00;
			16'hc75c: y = 16'hfe00;
			16'hc75d: y = 16'hfe00;
			16'hc75e: y = 16'hfe00;
			16'hc75f: y = 16'hfe00;
			16'hc760: y = 16'hfe00;
			16'hc761: y = 16'hfe00;
			16'hc762: y = 16'hfe00;
			16'hc763: y = 16'hfe00;
			16'hc764: y = 16'hfe00;
			16'hc765: y = 16'hfe00;
			16'hc766: y = 16'hfe00;
			16'hc767: y = 16'hfe00;
			16'hc768: y = 16'hfe00;
			16'hc769: y = 16'hfe00;
			16'hc76a: y = 16'hfe00;
			16'hc76b: y = 16'hfe00;
			16'hc76c: y = 16'hfe00;
			16'hc76d: y = 16'hfe00;
			16'hc76e: y = 16'hfe00;
			16'hc76f: y = 16'hfe00;
			16'hc770: y = 16'hfe00;
			16'hc771: y = 16'hfe00;
			16'hc772: y = 16'hfe00;
			16'hc773: y = 16'hfe00;
			16'hc774: y = 16'hfe00;
			16'hc775: y = 16'hfe00;
			16'hc776: y = 16'hfe00;
			16'hc777: y = 16'hfe00;
			16'hc778: y = 16'hfe00;
			16'hc779: y = 16'hfe00;
			16'hc77a: y = 16'hfe00;
			16'hc77b: y = 16'hfe00;
			16'hc77c: y = 16'hfe00;
			16'hc77d: y = 16'hfe00;
			16'hc77e: y = 16'hfe00;
			16'hc77f: y = 16'hfe00;
			16'hc780: y = 16'hfe00;
			16'hc781: y = 16'hfe00;
			16'hc782: y = 16'hfe00;
			16'hc783: y = 16'hfe00;
			16'hc784: y = 16'hfe00;
			16'hc785: y = 16'hfe00;
			16'hc786: y = 16'hfe00;
			16'hc787: y = 16'hfe00;
			16'hc788: y = 16'hfe00;
			16'hc789: y = 16'hfe00;
			16'hc78a: y = 16'hfe00;
			16'hc78b: y = 16'hfe00;
			16'hc78c: y = 16'hfe00;
			16'hc78d: y = 16'hfe00;
			16'hc78e: y = 16'hfe00;
			16'hc78f: y = 16'hfe00;
			16'hc790: y = 16'hfe00;
			16'hc791: y = 16'hfe00;
			16'hc792: y = 16'hfe00;
			16'hc793: y = 16'hfe00;
			16'hc794: y = 16'hfe00;
			16'hc795: y = 16'hfe00;
			16'hc796: y = 16'hfe00;
			16'hc797: y = 16'hfe00;
			16'hc798: y = 16'hfe00;
			16'hc799: y = 16'hfe00;
			16'hc79a: y = 16'hfe00;
			16'hc79b: y = 16'hfe00;
			16'hc79c: y = 16'hfe00;
			16'hc79d: y = 16'hfe00;
			16'hc79e: y = 16'hfe00;
			16'hc79f: y = 16'hfe00;
			16'hc7a0: y = 16'hfe00;
			16'hc7a1: y = 16'hfe00;
			16'hc7a2: y = 16'hfe00;
			16'hc7a3: y = 16'hfe00;
			16'hc7a4: y = 16'hfe00;
			16'hc7a5: y = 16'hfe00;
			16'hc7a6: y = 16'hfe00;
			16'hc7a7: y = 16'hfe00;
			16'hc7a8: y = 16'hfe00;
			16'hc7a9: y = 16'hfe00;
			16'hc7aa: y = 16'hfe00;
			16'hc7ab: y = 16'hfe00;
			16'hc7ac: y = 16'hfe00;
			16'hc7ad: y = 16'hfe00;
			16'hc7ae: y = 16'hfe00;
			16'hc7af: y = 16'hfe00;
			16'hc7b0: y = 16'hfe00;
			16'hc7b1: y = 16'hfe00;
			16'hc7b2: y = 16'hfe00;
			16'hc7b3: y = 16'hfe00;
			16'hc7b4: y = 16'hfe00;
			16'hc7b5: y = 16'hfe00;
			16'hc7b6: y = 16'hfe00;
			16'hc7b7: y = 16'hfe00;
			16'hc7b8: y = 16'hfe00;
			16'hc7b9: y = 16'hfe00;
			16'hc7ba: y = 16'hfe00;
			16'hc7bb: y = 16'hfe00;
			16'hc7bc: y = 16'hfe00;
			16'hc7bd: y = 16'hfe00;
			16'hc7be: y = 16'hfe00;
			16'hc7bf: y = 16'hfe00;
			16'hc7c0: y = 16'hfe00;
			16'hc7c1: y = 16'hfe00;
			16'hc7c2: y = 16'hfe00;
			16'hc7c3: y = 16'hfe00;
			16'hc7c4: y = 16'hfe00;
			16'hc7c5: y = 16'hfe00;
			16'hc7c6: y = 16'hfe00;
			16'hc7c7: y = 16'hfe00;
			16'hc7c8: y = 16'hfe00;
			16'hc7c9: y = 16'hfe00;
			16'hc7ca: y = 16'hfe00;
			16'hc7cb: y = 16'hfe00;
			16'hc7cc: y = 16'hfe00;
			16'hc7cd: y = 16'hfe00;
			16'hc7ce: y = 16'hfe00;
			16'hc7cf: y = 16'hfe00;
			16'hc7d0: y = 16'hfe00;
			16'hc7d1: y = 16'hfe00;
			16'hc7d2: y = 16'hfe00;
			16'hc7d3: y = 16'hfe00;
			16'hc7d4: y = 16'hfe00;
			16'hc7d5: y = 16'hfe00;
			16'hc7d6: y = 16'hfe00;
			16'hc7d7: y = 16'hfe00;
			16'hc7d8: y = 16'hfe00;
			16'hc7d9: y = 16'hfe00;
			16'hc7da: y = 16'hfe00;
			16'hc7db: y = 16'hfe00;
			16'hc7dc: y = 16'hfe00;
			16'hc7dd: y = 16'hfe00;
			16'hc7de: y = 16'hfe00;
			16'hc7df: y = 16'hfe00;
			16'hc7e0: y = 16'hfe00;
			16'hc7e1: y = 16'hfe00;
			16'hc7e2: y = 16'hfe00;
			16'hc7e3: y = 16'hfe00;
			16'hc7e4: y = 16'hfe00;
			16'hc7e5: y = 16'hfe00;
			16'hc7e6: y = 16'hfe00;
			16'hc7e7: y = 16'hfe00;
			16'hc7e8: y = 16'hfe00;
			16'hc7e9: y = 16'hfe00;
			16'hc7ea: y = 16'hfe00;
			16'hc7eb: y = 16'hfe00;
			16'hc7ec: y = 16'hfe00;
			16'hc7ed: y = 16'hfe00;
			16'hc7ee: y = 16'hfe00;
			16'hc7ef: y = 16'hfe00;
			16'hc7f0: y = 16'hfe00;
			16'hc7f1: y = 16'hfe00;
			16'hc7f2: y = 16'hfe00;
			16'hc7f3: y = 16'hfe00;
			16'hc7f4: y = 16'hfe00;
			16'hc7f5: y = 16'hfe00;
			16'hc7f6: y = 16'hfe00;
			16'hc7f7: y = 16'hfe00;
			16'hc7f8: y = 16'hfe00;
			16'hc7f9: y = 16'hfe00;
			16'hc7fa: y = 16'hfe00;
			16'hc7fb: y = 16'hfe00;
			16'hc7fc: y = 16'hfe00;
			16'hc7fd: y = 16'hfe00;
			16'hc7fe: y = 16'hfe00;
			16'hc7ff: y = 16'hfe00;
			16'hc800: y = 16'hfe00;
			16'hc801: y = 16'hfe00;
			16'hc802: y = 16'hfe00;
			16'hc803: y = 16'hfe00;
			16'hc804: y = 16'hfe00;
			16'hc805: y = 16'hfe00;
			16'hc806: y = 16'hfe00;
			16'hc807: y = 16'hfe00;
			16'hc808: y = 16'hfe00;
			16'hc809: y = 16'hfe00;
			16'hc80a: y = 16'hfe00;
			16'hc80b: y = 16'hfe00;
			16'hc80c: y = 16'hfe00;
			16'hc80d: y = 16'hfe00;
			16'hc80e: y = 16'hfe00;
			16'hc80f: y = 16'hfe00;
			16'hc810: y = 16'hfe00;
			16'hc811: y = 16'hfe00;
			16'hc812: y = 16'hfe00;
			16'hc813: y = 16'hfe00;
			16'hc814: y = 16'hfe00;
			16'hc815: y = 16'hfe00;
			16'hc816: y = 16'hfe00;
			16'hc817: y = 16'hfe00;
			16'hc818: y = 16'hfe00;
			16'hc819: y = 16'hfe00;
			16'hc81a: y = 16'hfe00;
			16'hc81b: y = 16'hfe00;
			16'hc81c: y = 16'hfe00;
			16'hc81d: y = 16'hfe00;
			16'hc81e: y = 16'hfe00;
			16'hc81f: y = 16'hfe00;
			16'hc820: y = 16'hfe00;
			16'hc821: y = 16'hfe00;
			16'hc822: y = 16'hfe00;
			16'hc823: y = 16'hfe00;
			16'hc824: y = 16'hfe00;
			16'hc825: y = 16'hfe00;
			16'hc826: y = 16'hfe00;
			16'hc827: y = 16'hfe00;
			16'hc828: y = 16'hfe00;
			16'hc829: y = 16'hfe00;
			16'hc82a: y = 16'hfe00;
			16'hc82b: y = 16'hfe00;
			16'hc82c: y = 16'hfe00;
			16'hc82d: y = 16'hfe00;
			16'hc82e: y = 16'hfe00;
			16'hc82f: y = 16'hfe00;
			16'hc830: y = 16'hfe00;
			16'hc831: y = 16'hfe00;
			16'hc832: y = 16'hfe00;
			16'hc833: y = 16'hfe00;
			16'hc834: y = 16'hfe00;
			16'hc835: y = 16'hfe00;
			16'hc836: y = 16'hfe00;
			16'hc837: y = 16'hfe00;
			16'hc838: y = 16'hfe00;
			16'hc839: y = 16'hfe00;
			16'hc83a: y = 16'hfe00;
			16'hc83b: y = 16'hfe00;
			16'hc83c: y = 16'hfe00;
			16'hc83d: y = 16'hfe00;
			16'hc83e: y = 16'hfe00;
			16'hc83f: y = 16'hfe00;
			16'hc840: y = 16'hfe00;
			16'hc841: y = 16'hfe00;
			16'hc842: y = 16'hfe00;
			16'hc843: y = 16'hfe00;
			16'hc844: y = 16'hfe00;
			16'hc845: y = 16'hfe00;
			16'hc846: y = 16'hfe00;
			16'hc847: y = 16'hfe00;
			16'hc848: y = 16'hfe00;
			16'hc849: y = 16'hfe00;
			16'hc84a: y = 16'hfe00;
			16'hc84b: y = 16'hfe00;
			16'hc84c: y = 16'hfe00;
			16'hc84d: y = 16'hfe00;
			16'hc84e: y = 16'hfe00;
			16'hc84f: y = 16'hfe00;
			16'hc850: y = 16'hfe00;
			16'hc851: y = 16'hfe00;
			16'hc852: y = 16'hfe00;
			16'hc853: y = 16'hfe00;
			16'hc854: y = 16'hfe00;
			16'hc855: y = 16'hfe00;
			16'hc856: y = 16'hfe00;
			16'hc857: y = 16'hfe00;
			16'hc858: y = 16'hfe00;
			16'hc859: y = 16'hfe00;
			16'hc85a: y = 16'hfe00;
			16'hc85b: y = 16'hfe00;
			16'hc85c: y = 16'hfe00;
			16'hc85d: y = 16'hfe00;
			16'hc85e: y = 16'hfe00;
			16'hc85f: y = 16'hfe00;
			16'hc860: y = 16'hfe00;
			16'hc861: y = 16'hfe00;
			16'hc862: y = 16'hfe00;
			16'hc863: y = 16'hfe00;
			16'hc864: y = 16'hfe00;
			16'hc865: y = 16'hfe00;
			16'hc866: y = 16'hfe00;
			16'hc867: y = 16'hfe00;
			16'hc868: y = 16'hfe00;
			16'hc869: y = 16'hfe00;
			16'hc86a: y = 16'hfe00;
			16'hc86b: y = 16'hfe00;
			16'hc86c: y = 16'hfe00;
			16'hc86d: y = 16'hfe00;
			16'hc86e: y = 16'hfe00;
			16'hc86f: y = 16'hfe00;
			16'hc870: y = 16'hfe00;
			16'hc871: y = 16'hfe00;
			16'hc872: y = 16'hfe00;
			16'hc873: y = 16'hfe00;
			16'hc874: y = 16'hfe00;
			16'hc875: y = 16'hfe00;
			16'hc876: y = 16'hfe00;
			16'hc877: y = 16'hfe00;
			16'hc878: y = 16'hfe00;
			16'hc879: y = 16'hfe00;
			16'hc87a: y = 16'hfe00;
			16'hc87b: y = 16'hfe00;
			16'hc87c: y = 16'hfe00;
			16'hc87d: y = 16'hfe00;
			16'hc87e: y = 16'hfe00;
			16'hc87f: y = 16'hfe00;
			16'hc880: y = 16'hfe00;
			16'hc881: y = 16'hfe00;
			16'hc882: y = 16'hfe00;
			16'hc883: y = 16'hfe00;
			16'hc884: y = 16'hfe00;
			16'hc885: y = 16'hfe00;
			16'hc886: y = 16'hfe00;
			16'hc887: y = 16'hfe00;
			16'hc888: y = 16'hfe00;
			16'hc889: y = 16'hfe00;
			16'hc88a: y = 16'hfe00;
			16'hc88b: y = 16'hfe00;
			16'hc88c: y = 16'hfe00;
			16'hc88d: y = 16'hfe00;
			16'hc88e: y = 16'hfe00;
			16'hc88f: y = 16'hfe00;
			16'hc890: y = 16'hfe00;
			16'hc891: y = 16'hfe00;
			16'hc892: y = 16'hfe00;
			16'hc893: y = 16'hfe00;
			16'hc894: y = 16'hfe00;
			16'hc895: y = 16'hfe00;
			16'hc896: y = 16'hfe00;
			16'hc897: y = 16'hfe00;
			16'hc898: y = 16'hfe00;
			16'hc899: y = 16'hfe00;
			16'hc89a: y = 16'hfe00;
			16'hc89b: y = 16'hfe00;
			16'hc89c: y = 16'hfe00;
			16'hc89d: y = 16'hfe00;
			16'hc89e: y = 16'hfe00;
			16'hc89f: y = 16'hfe00;
			16'hc8a0: y = 16'hfe00;
			16'hc8a1: y = 16'hfe00;
			16'hc8a2: y = 16'hfe00;
			16'hc8a3: y = 16'hfe00;
			16'hc8a4: y = 16'hfe00;
			16'hc8a5: y = 16'hfe00;
			16'hc8a6: y = 16'hfe00;
			16'hc8a7: y = 16'hfe00;
			16'hc8a8: y = 16'hfe00;
			16'hc8a9: y = 16'hfe00;
			16'hc8aa: y = 16'hfe00;
			16'hc8ab: y = 16'hfe00;
			16'hc8ac: y = 16'hfe00;
			16'hc8ad: y = 16'hfe00;
			16'hc8ae: y = 16'hfe00;
			16'hc8af: y = 16'hfe00;
			16'hc8b0: y = 16'hfe00;
			16'hc8b1: y = 16'hfe00;
			16'hc8b2: y = 16'hfe00;
			16'hc8b3: y = 16'hfe00;
			16'hc8b4: y = 16'hfe00;
			16'hc8b5: y = 16'hfe00;
			16'hc8b6: y = 16'hfe00;
			16'hc8b7: y = 16'hfe00;
			16'hc8b8: y = 16'hfe00;
			16'hc8b9: y = 16'hfe00;
			16'hc8ba: y = 16'hfe00;
			16'hc8bb: y = 16'hfe00;
			16'hc8bc: y = 16'hfe00;
			16'hc8bd: y = 16'hfe00;
			16'hc8be: y = 16'hfe00;
			16'hc8bf: y = 16'hfe00;
			16'hc8c0: y = 16'hfe00;
			16'hc8c1: y = 16'hfe00;
			16'hc8c2: y = 16'hfe00;
			16'hc8c3: y = 16'hfe00;
			16'hc8c4: y = 16'hfe00;
			16'hc8c5: y = 16'hfe00;
			16'hc8c6: y = 16'hfe00;
			16'hc8c7: y = 16'hfe00;
			16'hc8c8: y = 16'hfe00;
			16'hc8c9: y = 16'hfe00;
			16'hc8ca: y = 16'hfe00;
			16'hc8cb: y = 16'hfe00;
			16'hc8cc: y = 16'hfe00;
			16'hc8cd: y = 16'hfe00;
			16'hc8ce: y = 16'hfe00;
			16'hc8cf: y = 16'hfe00;
			16'hc8d0: y = 16'hfe00;
			16'hc8d1: y = 16'hfe00;
			16'hc8d2: y = 16'hfe00;
			16'hc8d3: y = 16'hfe00;
			16'hc8d4: y = 16'hfe00;
			16'hc8d5: y = 16'hfe00;
			16'hc8d6: y = 16'hfe00;
			16'hc8d7: y = 16'hfe00;
			16'hc8d8: y = 16'hfe00;
			16'hc8d9: y = 16'hfe00;
			16'hc8da: y = 16'hfe00;
			16'hc8db: y = 16'hfe00;
			16'hc8dc: y = 16'hfe00;
			16'hc8dd: y = 16'hfe00;
			16'hc8de: y = 16'hfe00;
			16'hc8df: y = 16'hfe00;
			16'hc8e0: y = 16'hfe00;
			16'hc8e1: y = 16'hfe00;
			16'hc8e2: y = 16'hfe00;
			16'hc8e3: y = 16'hfe00;
			16'hc8e4: y = 16'hfe00;
			16'hc8e5: y = 16'hfe00;
			16'hc8e6: y = 16'hfe00;
			16'hc8e7: y = 16'hfe00;
			16'hc8e8: y = 16'hfe00;
			16'hc8e9: y = 16'hfe00;
			16'hc8ea: y = 16'hfe00;
			16'hc8eb: y = 16'hfe00;
			16'hc8ec: y = 16'hfe00;
			16'hc8ed: y = 16'hfe00;
			16'hc8ee: y = 16'hfe00;
			16'hc8ef: y = 16'hfe00;
			16'hc8f0: y = 16'hfe00;
			16'hc8f1: y = 16'hfe00;
			16'hc8f2: y = 16'hfe00;
			16'hc8f3: y = 16'hfe00;
			16'hc8f4: y = 16'hfe00;
			16'hc8f5: y = 16'hfe00;
			16'hc8f6: y = 16'hfe00;
			16'hc8f7: y = 16'hfe00;
			16'hc8f8: y = 16'hfe00;
			16'hc8f9: y = 16'hfe00;
			16'hc8fa: y = 16'hfe00;
			16'hc8fb: y = 16'hfe00;
			16'hc8fc: y = 16'hfe00;
			16'hc8fd: y = 16'hfe00;
			16'hc8fe: y = 16'hfe00;
			16'hc8ff: y = 16'hfe00;
			16'hc900: y = 16'hfe00;
			16'hc901: y = 16'hfe00;
			16'hc902: y = 16'hfe00;
			16'hc903: y = 16'hfe00;
			16'hc904: y = 16'hfe00;
			16'hc905: y = 16'hfe00;
			16'hc906: y = 16'hfe00;
			16'hc907: y = 16'hfe00;
			16'hc908: y = 16'hfe00;
			16'hc909: y = 16'hfe00;
			16'hc90a: y = 16'hfe00;
			16'hc90b: y = 16'hfe00;
			16'hc90c: y = 16'hfe00;
			16'hc90d: y = 16'hfe00;
			16'hc90e: y = 16'hfe00;
			16'hc90f: y = 16'hfe00;
			16'hc910: y = 16'hfe00;
			16'hc911: y = 16'hfe00;
			16'hc912: y = 16'hfe00;
			16'hc913: y = 16'hfe00;
			16'hc914: y = 16'hfe00;
			16'hc915: y = 16'hfe00;
			16'hc916: y = 16'hfe00;
			16'hc917: y = 16'hfe00;
			16'hc918: y = 16'hfe00;
			16'hc919: y = 16'hfe00;
			16'hc91a: y = 16'hfe00;
			16'hc91b: y = 16'hfe00;
			16'hc91c: y = 16'hfe00;
			16'hc91d: y = 16'hfe00;
			16'hc91e: y = 16'hfe00;
			16'hc91f: y = 16'hfe00;
			16'hc920: y = 16'hfe00;
			16'hc921: y = 16'hfe00;
			16'hc922: y = 16'hfe00;
			16'hc923: y = 16'hfe00;
			16'hc924: y = 16'hfe00;
			16'hc925: y = 16'hfe00;
			16'hc926: y = 16'hfe00;
			16'hc927: y = 16'hfe00;
			16'hc928: y = 16'hfe00;
			16'hc929: y = 16'hfe00;
			16'hc92a: y = 16'hfe00;
			16'hc92b: y = 16'hfe00;
			16'hc92c: y = 16'hfe00;
			16'hc92d: y = 16'hfe00;
			16'hc92e: y = 16'hfe00;
			16'hc92f: y = 16'hfe00;
			16'hc930: y = 16'hfe00;
			16'hc931: y = 16'hfe00;
			16'hc932: y = 16'hfe00;
			16'hc933: y = 16'hfe00;
			16'hc934: y = 16'hfe00;
			16'hc935: y = 16'hfe00;
			16'hc936: y = 16'hfe00;
			16'hc937: y = 16'hfe00;
			16'hc938: y = 16'hfe00;
			16'hc939: y = 16'hfe00;
			16'hc93a: y = 16'hfe00;
			16'hc93b: y = 16'hfe00;
			16'hc93c: y = 16'hfe00;
			16'hc93d: y = 16'hfe00;
			16'hc93e: y = 16'hfe00;
			16'hc93f: y = 16'hfe00;
			16'hc940: y = 16'hfe00;
			16'hc941: y = 16'hfe00;
			16'hc942: y = 16'hfe00;
			16'hc943: y = 16'hfe00;
			16'hc944: y = 16'hfe00;
			16'hc945: y = 16'hfe00;
			16'hc946: y = 16'hfe00;
			16'hc947: y = 16'hfe00;
			16'hc948: y = 16'hfe00;
			16'hc949: y = 16'hfe00;
			16'hc94a: y = 16'hfe00;
			16'hc94b: y = 16'hfe00;
			16'hc94c: y = 16'hfe00;
			16'hc94d: y = 16'hfe00;
			16'hc94e: y = 16'hfe00;
			16'hc94f: y = 16'hfe00;
			16'hc950: y = 16'hfe00;
			16'hc951: y = 16'hfe00;
			16'hc952: y = 16'hfe00;
			16'hc953: y = 16'hfe00;
			16'hc954: y = 16'hfe00;
			16'hc955: y = 16'hfe00;
			16'hc956: y = 16'hfe00;
			16'hc957: y = 16'hfe00;
			16'hc958: y = 16'hfe00;
			16'hc959: y = 16'hfe00;
			16'hc95a: y = 16'hfe00;
			16'hc95b: y = 16'hfe00;
			16'hc95c: y = 16'hfe00;
			16'hc95d: y = 16'hfe00;
			16'hc95e: y = 16'hfe00;
			16'hc95f: y = 16'hfe00;
			16'hc960: y = 16'hfe00;
			16'hc961: y = 16'hfe00;
			16'hc962: y = 16'hfe00;
			16'hc963: y = 16'hfe00;
			16'hc964: y = 16'hfe00;
			16'hc965: y = 16'hfe00;
			16'hc966: y = 16'hfe00;
			16'hc967: y = 16'hfe00;
			16'hc968: y = 16'hfe00;
			16'hc969: y = 16'hfe00;
			16'hc96a: y = 16'hfe00;
			16'hc96b: y = 16'hfe00;
			16'hc96c: y = 16'hfe00;
			16'hc96d: y = 16'hfe00;
			16'hc96e: y = 16'hfe00;
			16'hc96f: y = 16'hfe00;
			16'hc970: y = 16'hfe00;
			16'hc971: y = 16'hfe00;
			16'hc972: y = 16'hfe00;
			16'hc973: y = 16'hfe00;
			16'hc974: y = 16'hfe00;
			16'hc975: y = 16'hfe00;
			16'hc976: y = 16'hfe00;
			16'hc977: y = 16'hfe00;
			16'hc978: y = 16'hfe00;
			16'hc979: y = 16'hfe00;
			16'hc97a: y = 16'hfe00;
			16'hc97b: y = 16'hfe00;
			16'hc97c: y = 16'hfe00;
			16'hc97d: y = 16'hfe00;
			16'hc97e: y = 16'hfe00;
			16'hc97f: y = 16'hfe00;
			16'hc980: y = 16'hfe00;
			16'hc981: y = 16'hfe00;
			16'hc982: y = 16'hfe00;
			16'hc983: y = 16'hfe00;
			16'hc984: y = 16'hfe00;
			16'hc985: y = 16'hfe00;
			16'hc986: y = 16'hfe00;
			16'hc987: y = 16'hfe00;
			16'hc988: y = 16'hfe00;
			16'hc989: y = 16'hfe00;
			16'hc98a: y = 16'hfe00;
			16'hc98b: y = 16'hfe00;
			16'hc98c: y = 16'hfe00;
			16'hc98d: y = 16'hfe00;
			16'hc98e: y = 16'hfe00;
			16'hc98f: y = 16'hfe00;
			16'hc990: y = 16'hfe00;
			16'hc991: y = 16'hfe00;
			16'hc992: y = 16'hfe00;
			16'hc993: y = 16'hfe00;
			16'hc994: y = 16'hfe00;
			16'hc995: y = 16'hfe00;
			16'hc996: y = 16'hfe00;
			16'hc997: y = 16'hfe00;
			16'hc998: y = 16'hfe00;
			16'hc999: y = 16'hfe00;
			16'hc99a: y = 16'hfe00;
			16'hc99b: y = 16'hfe00;
			16'hc99c: y = 16'hfe00;
			16'hc99d: y = 16'hfe00;
			16'hc99e: y = 16'hfe00;
			16'hc99f: y = 16'hfe00;
			16'hc9a0: y = 16'hfe00;
			16'hc9a1: y = 16'hfe00;
			16'hc9a2: y = 16'hfe00;
			16'hc9a3: y = 16'hfe00;
			16'hc9a4: y = 16'hfe00;
			16'hc9a5: y = 16'hfe00;
			16'hc9a6: y = 16'hfe00;
			16'hc9a7: y = 16'hfe00;
			16'hc9a8: y = 16'hfe00;
			16'hc9a9: y = 16'hfe00;
			16'hc9aa: y = 16'hfe00;
			16'hc9ab: y = 16'hfe00;
			16'hc9ac: y = 16'hfe00;
			16'hc9ad: y = 16'hfe00;
			16'hc9ae: y = 16'hfe00;
			16'hc9af: y = 16'hfe00;
			16'hc9b0: y = 16'hfe00;
			16'hc9b1: y = 16'hfe00;
			16'hc9b2: y = 16'hfe00;
			16'hc9b3: y = 16'hfe00;
			16'hc9b4: y = 16'hfe00;
			16'hc9b5: y = 16'hfe00;
			16'hc9b6: y = 16'hfe00;
			16'hc9b7: y = 16'hfe00;
			16'hc9b8: y = 16'hfe00;
			16'hc9b9: y = 16'hfe00;
			16'hc9ba: y = 16'hfe00;
			16'hc9bb: y = 16'hfe00;
			16'hc9bc: y = 16'hfe00;
			16'hc9bd: y = 16'hfe00;
			16'hc9be: y = 16'hfe00;
			16'hc9bf: y = 16'hfe00;
			16'hc9c0: y = 16'hfe00;
			16'hc9c1: y = 16'hfe00;
			16'hc9c2: y = 16'hfe00;
			16'hc9c3: y = 16'hfe00;
			16'hc9c4: y = 16'hfe00;
			16'hc9c5: y = 16'hfe00;
			16'hc9c6: y = 16'hfe00;
			16'hc9c7: y = 16'hfe00;
			16'hc9c8: y = 16'hfe00;
			16'hc9c9: y = 16'hfe00;
			16'hc9ca: y = 16'hfe00;
			16'hc9cb: y = 16'hfe00;
			16'hc9cc: y = 16'hfe00;
			16'hc9cd: y = 16'hfe00;
			16'hc9ce: y = 16'hfe00;
			16'hc9cf: y = 16'hfe00;
			16'hc9d0: y = 16'hfe00;
			16'hc9d1: y = 16'hfe00;
			16'hc9d2: y = 16'hfe00;
			16'hc9d3: y = 16'hfe00;
			16'hc9d4: y = 16'hfe00;
			16'hc9d5: y = 16'hfe00;
			16'hc9d6: y = 16'hfe00;
			16'hc9d7: y = 16'hfe00;
			16'hc9d8: y = 16'hfe00;
			16'hc9d9: y = 16'hfe00;
			16'hc9da: y = 16'hfe00;
			16'hc9db: y = 16'hfe00;
			16'hc9dc: y = 16'hfe00;
			16'hc9dd: y = 16'hfe00;
			16'hc9de: y = 16'hfe00;
			16'hc9df: y = 16'hfe00;
			16'hc9e0: y = 16'hfe00;
			16'hc9e1: y = 16'hfe00;
			16'hc9e2: y = 16'hfe00;
			16'hc9e3: y = 16'hfe00;
			16'hc9e4: y = 16'hfe00;
			16'hc9e5: y = 16'hfe00;
			16'hc9e6: y = 16'hfe00;
			16'hc9e7: y = 16'hfe00;
			16'hc9e8: y = 16'hfe00;
			16'hc9e9: y = 16'hfe00;
			16'hc9ea: y = 16'hfe00;
			16'hc9eb: y = 16'hfe00;
			16'hc9ec: y = 16'hfe00;
			16'hc9ed: y = 16'hfe00;
			16'hc9ee: y = 16'hfe00;
			16'hc9ef: y = 16'hfe00;
			16'hc9f0: y = 16'hfe00;
			16'hc9f1: y = 16'hfe00;
			16'hc9f2: y = 16'hfe00;
			16'hc9f3: y = 16'hfe00;
			16'hc9f4: y = 16'hfe00;
			16'hc9f5: y = 16'hfe00;
			16'hc9f6: y = 16'hfe00;
			16'hc9f7: y = 16'hfe00;
			16'hc9f8: y = 16'hfe00;
			16'hc9f9: y = 16'hfe00;
			16'hc9fa: y = 16'hfe00;
			16'hc9fb: y = 16'hfe00;
			16'hc9fc: y = 16'hfe00;
			16'hc9fd: y = 16'hfe00;
			16'hc9fe: y = 16'hfe00;
			16'hc9ff: y = 16'hfe00;
			16'hca00: y = 16'hfe00;
			16'hca01: y = 16'hfe00;
			16'hca02: y = 16'hfe00;
			16'hca03: y = 16'hfe00;
			16'hca04: y = 16'hfe00;
			16'hca05: y = 16'hfe00;
			16'hca06: y = 16'hfe00;
			16'hca07: y = 16'hfe00;
			16'hca08: y = 16'hfe00;
			16'hca09: y = 16'hfe00;
			16'hca0a: y = 16'hfe00;
			16'hca0b: y = 16'hfe00;
			16'hca0c: y = 16'hfe00;
			16'hca0d: y = 16'hfe00;
			16'hca0e: y = 16'hfe00;
			16'hca0f: y = 16'hfe00;
			16'hca10: y = 16'hfe00;
			16'hca11: y = 16'hfe00;
			16'hca12: y = 16'hfe00;
			16'hca13: y = 16'hfe00;
			16'hca14: y = 16'hfe00;
			16'hca15: y = 16'hfe00;
			16'hca16: y = 16'hfe00;
			16'hca17: y = 16'hfe00;
			16'hca18: y = 16'hfe00;
			16'hca19: y = 16'hfe00;
			16'hca1a: y = 16'hfe00;
			16'hca1b: y = 16'hfe00;
			16'hca1c: y = 16'hfe00;
			16'hca1d: y = 16'hfe00;
			16'hca1e: y = 16'hfe00;
			16'hca1f: y = 16'hfe00;
			16'hca20: y = 16'hfe00;
			16'hca21: y = 16'hfe00;
			16'hca22: y = 16'hfe00;
			16'hca23: y = 16'hfe00;
			16'hca24: y = 16'hfe00;
			16'hca25: y = 16'hfe00;
			16'hca26: y = 16'hfe00;
			16'hca27: y = 16'hfe00;
			16'hca28: y = 16'hfe00;
			16'hca29: y = 16'hfe00;
			16'hca2a: y = 16'hfe00;
			16'hca2b: y = 16'hfe00;
			16'hca2c: y = 16'hfe00;
			16'hca2d: y = 16'hfe00;
			16'hca2e: y = 16'hfe00;
			16'hca2f: y = 16'hfe00;
			16'hca30: y = 16'hfe00;
			16'hca31: y = 16'hfe00;
			16'hca32: y = 16'hfe00;
			16'hca33: y = 16'hfe00;
			16'hca34: y = 16'hfe00;
			16'hca35: y = 16'hfe00;
			16'hca36: y = 16'hfe00;
			16'hca37: y = 16'hfe00;
			16'hca38: y = 16'hfe00;
			16'hca39: y = 16'hfe00;
			16'hca3a: y = 16'hfe00;
			16'hca3b: y = 16'hfe00;
			16'hca3c: y = 16'hfe00;
			16'hca3d: y = 16'hfe00;
			16'hca3e: y = 16'hfe00;
			16'hca3f: y = 16'hfe00;
			16'hca40: y = 16'hfe00;
			16'hca41: y = 16'hfe00;
			16'hca42: y = 16'hfe00;
			16'hca43: y = 16'hfe00;
			16'hca44: y = 16'hfe00;
			16'hca45: y = 16'hfe00;
			16'hca46: y = 16'hfe00;
			16'hca47: y = 16'hfe00;
			16'hca48: y = 16'hfe00;
			16'hca49: y = 16'hfe00;
			16'hca4a: y = 16'hfe00;
			16'hca4b: y = 16'hfe00;
			16'hca4c: y = 16'hfe00;
			16'hca4d: y = 16'hfe00;
			16'hca4e: y = 16'hfe00;
			16'hca4f: y = 16'hfe00;
			16'hca50: y = 16'hfe00;
			16'hca51: y = 16'hfe00;
			16'hca52: y = 16'hfe00;
			16'hca53: y = 16'hfe00;
			16'hca54: y = 16'hfe00;
			16'hca55: y = 16'hfe00;
			16'hca56: y = 16'hfe00;
			16'hca57: y = 16'hfe00;
			16'hca58: y = 16'hfe00;
			16'hca59: y = 16'hfe00;
			16'hca5a: y = 16'hfe00;
			16'hca5b: y = 16'hfe00;
			16'hca5c: y = 16'hfe00;
			16'hca5d: y = 16'hfe00;
			16'hca5e: y = 16'hfe00;
			16'hca5f: y = 16'hfe00;
			16'hca60: y = 16'hfe00;
			16'hca61: y = 16'hfe00;
			16'hca62: y = 16'hfe00;
			16'hca63: y = 16'hfe00;
			16'hca64: y = 16'hfe00;
			16'hca65: y = 16'hfe00;
			16'hca66: y = 16'hfe00;
			16'hca67: y = 16'hfe00;
			16'hca68: y = 16'hfe00;
			16'hca69: y = 16'hfe00;
			16'hca6a: y = 16'hfe00;
			16'hca6b: y = 16'hfe00;
			16'hca6c: y = 16'hfe00;
			16'hca6d: y = 16'hfe00;
			16'hca6e: y = 16'hfe00;
			16'hca6f: y = 16'hfe00;
			16'hca70: y = 16'hfe00;
			16'hca71: y = 16'hfe00;
			16'hca72: y = 16'hfe00;
			16'hca73: y = 16'hfe00;
			16'hca74: y = 16'hfe00;
			16'hca75: y = 16'hfe00;
			16'hca76: y = 16'hfe00;
			16'hca77: y = 16'hfe00;
			16'hca78: y = 16'hfe00;
			16'hca79: y = 16'hfe00;
			16'hca7a: y = 16'hfe00;
			16'hca7b: y = 16'hfe00;
			16'hca7c: y = 16'hfe00;
			16'hca7d: y = 16'hfe00;
			16'hca7e: y = 16'hfe00;
			16'hca7f: y = 16'hfe00;
			16'hca80: y = 16'hfe00;
			16'hca81: y = 16'hfe00;
			16'hca82: y = 16'hfe00;
			16'hca83: y = 16'hfe00;
			16'hca84: y = 16'hfe00;
			16'hca85: y = 16'hfe00;
			16'hca86: y = 16'hfe00;
			16'hca87: y = 16'hfe00;
			16'hca88: y = 16'hfe00;
			16'hca89: y = 16'hfe00;
			16'hca8a: y = 16'hfe00;
			16'hca8b: y = 16'hfe00;
			16'hca8c: y = 16'hfe00;
			16'hca8d: y = 16'hfe00;
			16'hca8e: y = 16'hfe00;
			16'hca8f: y = 16'hfe00;
			16'hca90: y = 16'hfe00;
			16'hca91: y = 16'hfe00;
			16'hca92: y = 16'hfe00;
			16'hca93: y = 16'hfe00;
			16'hca94: y = 16'hfe00;
			16'hca95: y = 16'hfe00;
			16'hca96: y = 16'hfe00;
			16'hca97: y = 16'hfe00;
			16'hca98: y = 16'hfe00;
			16'hca99: y = 16'hfe00;
			16'hca9a: y = 16'hfe00;
			16'hca9b: y = 16'hfe00;
			16'hca9c: y = 16'hfe00;
			16'hca9d: y = 16'hfe00;
			16'hca9e: y = 16'hfe00;
			16'hca9f: y = 16'hfe00;
			16'hcaa0: y = 16'hfe00;
			16'hcaa1: y = 16'hfe00;
			16'hcaa2: y = 16'hfe00;
			16'hcaa3: y = 16'hfe00;
			16'hcaa4: y = 16'hfe00;
			16'hcaa5: y = 16'hfe00;
			16'hcaa6: y = 16'hfe00;
			16'hcaa7: y = 16'hfe00;
			16'hcaa8: y = 16'hfe00;
			16'hcaa9: y = 16'hfe00;
			16'hcaaa: y = 16'hfe00;
			16'hcaab: y = 16'hfe00;
			16'hcaac: y = 16'hfe00;
			16'hcaad: y = 16'hfe00;
			16'hcaae: y = 16'hfe00;
			16'hcaaf: y = 16'hfe00;
			16'hcab0: y = 16'hfe00;
			16'hcab1: y = 16'hfe00;
			16'hcab2: y = 16'hfe00;
			16'hcab3: y = 16'hfe00;
			16'hcab4: y = 16'hfe00;
			16'hcab5: y = 16'hfe00;
			16'hcab6: y = 16'hfe00;
			16'hcab7: y = 16'hfe00;
			16'hcab8: y = 16'hfe00;
			16'hcab9: y = 16'hfe00;
			16'hcaba: y = 16'hfe00;
			16'hcabb: y = 16'hfe00;
			16'hcabc: y = 16'hfe00;
			16'hcabd: y = 16'hfe00;
			16'hcabe: y = 16'hfe00;
			16'hcabf: y = 16'hfe00;
			16'hcac0: y = 16'hfe00;
			16'hcac1: y = 16'hfe00;
			16'hcac2: y = 16'hfe00;
			16'hcac3: y = 16'hfe00;
			16'hcac4: y = 16'hfe00;
			16'hcac5: y = 16'hfe00;
			16'hcac6: y = 16'hfe00;
			16'hcac7: y = 16'hfe00;
			16'hcac8: y = 16'hfe00;
			16'hcac9: y = 16'hfe00;
			16'hcaca: y = 16'hfe00;
			16'hcacb: y = 16'hfe00;
			16'hcacc: y = 16'hfe00;
			16'hcacd: y = 16'hfe00;
			16'hcace: y = 16'hfe00;
			16'hcacf: y = 16'hfe00;
			16'hcad0: y = 16'hfe00;
			16'hcad1: y = 16'hfe00;
			16'hcad2: y = 16'hfe00;
			16'hcad3: y = 16'hfe00;
			16'hcad4: y = 16'hfe00;
			16'hcad5: y = 16'hfe00;
			16'hcad6: y = 16'hfe00;
			16'hcad7: y = 16'hfe00;
			16'hcad8: y = 16'hfe00;
			16'hcad9: y = 16'hfe00;
			16'hcada: y = 16'hfe00;
			16'hcadb: y = 16'hfe00;
			16'hcadc: y = 16'hfe00;
			16'hcadd: y = 16'hfe00;
			16'hcade: y = 16'hfe00;
			16'hcadf: y = 16'hfe00;
			16'hcae0: y = 16'hfe00;
			16'hcae1: y = 16'hfe00;
			16'hcae2: y = 16'hfe00;
			16'hcae3: y = 16'hfe00;
			16'hcae4: y = 16'hfe00;
			16'hcae5: y = 16'hfe00;
			16'hcae6: y = 16'hfe00;
			16'hcae7: y = 16'hfe00;
			16'hcae8: y = 16'hfe00;
			16'hcae9: y = 16'hfe00;
			16'hcaea: y = 16'hfe00;
			16'hcaeb: y = 16'hfe00;
			16'hcaec: y = 16'hfe00;
			16'hcaed: y = 16'hfe00;
			16'hcaee: y = 16'hfe00;
			16'hcaef: y = 16'hfe00;
			16'hcaf0: y = 16'hfe00;
			16'hcaf1: y = 16'hfe00;
			16'hcaf2: y = 16'hfe00;
			16'hcaf3: y = 16'hfe00;
			16'hcaf4: y = 16'hfe00;
			16'hcaf5: y = 16'hfe00;
			16'hcaf6: y = 16'hfe00;
			16'hcaf7: y = 16'hfe00;
			16'hcaf8: y = 16'hfe00;
			16'hcaf9: y = 16'hfe00;
			16'hcafa: y = 16'hfe00;
			16'hcafb: y = 16'hfe00;
			16'hcafc: y = 16'hfe00;
			16'hcafd: y = 16'hfe00;
			16'hcafe: y = 16'hfe00;
			16'hcaff: y = 16'hfe00;
			16'hcb00: y = 16'hfe00;
			16'hcb01: y = 16'hfe00;
			16'hcb02: y = 16'hfe00;
			16'hcb03: y = 16'hfe00;
			16'hcb04: y = 16'hfe00;
			16'hcb05: y = 16'hfe00;
			16'hcb06: y = 16'hfe00;
			16'hcb07: y = 16'hfe00;
			16'hcb08: y = 16'hfe00;
			16'hcb09: y = 16'hfe00;
			16'hcb0a: y = 16'hfe00;
			16'hcb0b: y = 16'hfe00;
			16'hcb0c: y = 16'hfe00;
			16'hcb0d: y = 16'hfe00;
			16'hcb0e: y = 16'hfe00;
			16'hcb0f: y = 16'hfe00;
			16'hcb10: y = 16'hfe00;
			16'hcb11: y = 16'hfe00;
			16'hcb12: y = 16'hfe00;
			16'hcb13: y = 16'hfe00;
			16'hcb14: y = 16'hfe00;
			16'hcb15: y = 16'hfe00;
			16'hcb16: y = 16'hfe00;
			16'hcb17: y = 16'hfe00;
			16'hcb18: y = 16'hfe00;
			16'hcb19: y = 16'hfe00;
			16'hcb1a: y = 16'hfe00;
			16'hcb1b: y = 16'hfe00;
			16'hcb1c: y = 16'hfe00;
			16'hcb1d: y = 16'hfe00;
			16'hcb1e: y = 16'hfe00;
			16'hcb1f: y = 16'hfe00;
			16'hcb20: y = 16'hfe00;
			16'hcb21: y = 16'hfe00;
			16'hcb22: y = 16'hfe00;
			16'hcb23: y = 16'hfe00;
			16'hcb24: y = 16'hfe00;
			16'hcb25: y = 16'hfe00;
			16'hcb26: y = 16'hfe00;
			16'hcb27: y = 16'hfe00;
			16'hcb28: y = 16'hfe00;
			16'hcb29: y = 16'hfe00;
			16'hcb2a: y = 16'hfe00;
			16'hcb2b: y = 16'hfe00;
			16'hcb2c: y = 16'hfe00;
			16'hcb2d: y = 16'hfe00;
			16'hcb2e: y = 16'hfe00;
			16'hcb2f: y = 16'hfe00;
			16'hcb30: y = 16'hfe00;
			16'hcb31: y = 16'hfe00;
			16'hcb32: y = 16'hfe00;
			16'hcb33: y = 16'hfe00;
			16'hcb34: y = 16'hfe00;
			16'hcb35: y = 16'hfe00;
			16'hcb36: y = 16'hfe00;
			16'hcb37: y = 16'hfe00;
			16'hcb38: y = 16'hfe00;
			16'hcb39: y = 16'hfe00;
			16'hcb3a: y = 16'hfe00;
			16'hcb3b: y = 16'hfe00;
			16'hcb3c: y = 16'hfe00;
			16'hcb3d: y = 16'hfe00;
			16'hcb3e: y = 16'hfe00;
			16'hcb3f: y = 16'hfe00;
			16'hcb40: y = 16'hfe00;
			16'hcb41: y = 16'hfe00;
			16'hcb42: y = 16'hfe00;
			16'hcb43: y = 16'hfe00;
			16'hcb44: y = 16'hfe00;
			16'hcb45: y = 16'hfe00;
			16'hcb46: y = 16'hfe00;
			16'hcb47: y = 16'hfe00;
			16'hcb48: y = 16'hfe00;
			16'hcb49: y = 16'hfe00;
			16'hcb4a: y = 16'hfe00;
			16'hcb4b: y = 16'hfe00;
			16'hcb4c: y = 16'hfe00;
			16'hcb4d: y = 16'hfe00;
			16'hcb4e: y = 16'hfe00;
			16'hcb4f: y = 16'hfe00;
			16'hcb50: y = 16'hfe00;
			16'hcb51: y = 16'hfe00;
			16'hcb52: y = 16'hfe00;
			16'hcb53: y = 16'hfe00;
			16'hcb54: y = 16'hfe00;
			16'hcb55: y = 16'hfe00;
			16'hcb56: y = 16'hfe00;
			16'hcb57: y = 16'hfe00;
			16'hcb58: y = 16'hfe00;
			16'hcb59: y = 16'hfe00;
			16'hcb5a: y = 16'hfe00;
			16'hcb5b: y = 16'hfe00;
			16'hcb5c: y = 16'hfe00;
			16'hcb5d: y = 16'hfe00;
			16'hcb5e: y = 16'hfe00;
			16'hcb5f: y = 16'hfe00;
			16'hcb60: y = 16'hfe00;
			16'hcb61: y = 16'hfe00;
			16'hcb62: y = 16'hfe00;
			16'hcb63: y = 16'hfe00;
			16'hcb64: y = 16'hfe00;
			16'hcb65: y = 16'hfe00;
			16'hcb66: y = 16'hfe00;
			16'hcb67: y = 16'hfe00;
			16'hcb68: y = 16'hfe00;
			16'hcb69: y = 16'hfe00;
			16'hcb6a: y = 16'hfe00;
			16'hcb6b: y = 16'hfe00;
			16'hcb6c: y = 16'hfe00;
			16'hcb6d: y = 16'hfe00;
			16'hcb6e: y = 16'hfe00;
			16'hcb6f: y = 16'hfe00;
			16'hcb70: y = 16'hfe00;
			16'hcb71: y = 16'hfe00;
			16'hcb72: y = 16'hfe00;
			16'hcb73: y = 16'hfe00;
			16'hcb74: y = 16'hfe00;
			16'hcb75: y = 16'hfe00;
			16'hcb76: y = 16'hfe00;
			16'hcb77: y = 16'hfe00;
			16'hcb78: y = 16'hfe00;
			16'hcb79: y = 16'hfe00;
			16'hcb7a: y = 16'hfe00;
			16'hcb7b: y = 16'hfe00;
			16'hcb7c: y = 16'hfe00;
			16'hcb7d: y = 16'hfe00;
			16'hcb7e: y = 16'hfe00;
			16'hcb7f: y = 16'hfe00;
			16'hcb80: y = 16'hfe00;
			16'hcb81: y = 16'hfe00;
			16'hcb82: y = 16'hfe00;
			16'hcb83: y = 16'hfe00;
			16'hcb84: y = 16'hfe00;
			16'hcb85: y = 16'hfe00;
			16'hcb86: y = 16'hfe00;
			16'hcb87: y = 16'hfe00;
			16'hcb88: y = 16'hfe00;
			16'hcb89: y = 16'hfe00;
			16'hcb8a: y = 16'hfe00;
			16'hcb8b: y = 16'hfe00;
			16'hcb8c: y = 16'hfe00;
			16'hcb8d: y = 16'hfe00;
			16'hcb8e: y = 16'hfe00;
			16'hcb8f: y = 16'hfe00;
			16'hcb90: y = 16'hfe00;
			16'hcb91: y = 16'hfe00;
			16'hcb92: y = 16'hfe00;
			16'hcb93: y = 16'hfe00;
			16'hcb94: y = 16'hfe00;
			16'hcb95: y = 16'hfe00;
			16'hcb96: y = 16'hfe00;
			16'hcb97: y = 16'hfe00;
			16'hcb98: y = 16'hfe00;
			16'hcb99: y = 16'hfe00;
			16'hcb9a: y = 16'hfe00;
			16'hcb9b: y = 16'hfe00;
			16'hcb9c: y = 16'hfe00;
			16'hcb9d: y = 16'hfe00;
			16'hcb9e: y = 16'hfe00;
			16'hcb9f: y = 16'hfe00;
			16'hcba0: y = 16'hfe00;
			16'hcba1: y = 16'hfe00;
			16'hcba2: y = 16'hfe00;
			16'hcba3: y = 16'hfe00;
			16'hcba4: y = 16'hfe00;
			16'hcba5: y = 16'hfe00;
			16'hcba6: y = 16'hfe00;
			16'hcba7: y = 16'hfe00;
			16'hcba8: y = 16'hfe00;
			16'hcba9: y = 16'hfe00;
			16'hcbaa: y = 16'hfe00;
			16'hcbab: y = 16'hfe00;
			16'hcbac: y = 16'hfe00;
			16'hcbad: y = 16'hfe00;
			16'hcbae: y = 16'hfe00;
			16'hcbaf: y = 16'hfe00;
			16'hcbb0: y = 16'hfe00;
			16'hcbb1: y = 16'hfe00;
			16'hcbb2: y = 16'hfe00;
			16'hcbb3: y = 16'hfe00;
			16'hcbb4: y = 16'hfe00;
			16'hcbb5: y = 16'hfe00;
			16'hcbb6: y = 16'hfe00;
			16'hcbb7: y = 16'hfe00;
			16'hcbb8: y = 16'hfe00;
			16'hcbb9: y = 16'hfe00;
			16'hcbba: y = 16'hfe00;
			16'hcbbb: y = 16'hfe00;
			16'hcbbc: y = 16'hfe00;
			16'hcbbd: y = 16'hfe00;
			16'hcbbe: y = 16'hfe00;
			16'hcbbf: y = 16'hfe00;
			16'hcbc0: y = 16'hfe00;
			16'hcbc1: y = 16'hfe00;
			16'hcbc2: y = 16'hfe00;
			16'hcbc3: y = 16'hfe00;
			16'hcbc4: y = 16'hfe00;
			16'hcbc5: y = 16'hfe00;
			16'hcbc6: y = 16'hfe00;
			16'hcbc7: y = 16'hfe00;
			16'hcbc8: y = 16'hfe00;
			16'hcbc9: y = 16'hfe00;
			16'hcbca: y = 16'hfe00;
			16'hcbcb: y = 16'hfe00;
			16'hcbcc: y = 16'hfe00;
			16'hcbcd: y = 16'hfe00;
			16'hcbce: y = 16'hfe00;
			16'hcbcf: y = 16'hfe00;
			16'hcbd0: y = 16'hfe00;
			16'hcbd1: y = 16'hfe00;
			16'hcbd2: y = 16'hfe00;
			16'hcbd3: y = 16'hfe00;
			16'hcbd4: y = 16'hfe00;
			16'hcbd5: y = 16'hfe00;
			16'hcbd6: y = 16'hfe00;
			16'hcbd7: y = 16'hfe00;
			16'hcbd8: y = 16'hfe00;
			16'hcbd9: y = 16'hfe00;
			16'hcbda: y = 16'hfe00;
			16'hcbdb: y = 16'hfe00;
			16'hcbdc: y = 16'hfe00;
			16'hcbdd: y = 16'hfe00;
			16'hcbde: y = 16'hfe00;
			16'hcbdf: y = 16'hfe00;
			16'hcbe0: y = 16'hfe00;
			16'hcbe1: y = 16'hfe00;
			16'hcbe2: y = 16'hfe00;
			16'hcbe3: y = 16'hfe00;
			16'hcbe4: y = 16'hfe00;
			16'hcbe5: y = 16'hfe00;
			16'hcbe6: y = 16'hfe00;
			16'hcbe7: y = 16'hfe00;
			16'hcbe8: y = 16'hfe00;
			16'hcbe9: y = 16'hfe00;
			16'hcbea: y = 16'hfe00;
			16'hcbeb: y = 16'hfe00;
			16'hcbec: y = 16'hfe00;
			16'hcbed: y = 16'hfe00;
			16'hcbee: y = 16'hfe00;
			16'hcbef: y = 16'hfe00;
			16'hcbf0: y = 16'hfe00;
			16'hcbf1: y = 16'hfe00;
			16'hcbf2: y = 16'hfe00;
			16'hcbf3: y = 16'hfe00;
			16'hcbf4: y = 16'hfe00;
			16'hcbf5: y = 16'hfe00;
			16'hcbf6: y = 16'hfe00;
			16'hcbf7: y = 16'hfe00;
			16'hcbf8: y = 16'hfe00;
			16'hcbf9: y = 16'hfe00;
			16'hcbfa: y = 16'hfe00;
			16'hcbfb: y = 16'hfe00;
			16'hcbfc: y = 16'hfe00;
			16'hcbfd: y = 16'hfe00;
			16'hcbfe: y = 16'hfe00;
			16'hcbff: y = 16'hfe00;
			16'hcc00: y = 16'hfe00;
			16'hcc01: y = 16'hfe00;
			16'hcc02: y = 16'hfe00;
			16'hcc03: y = 16'hfe00;
			16'hcc04: y = 16'hfe00;
			16'hcc05: y = 16'hfe00;
			16'hcc06: y = 16'hfe00;
			16'hcc07: y = 16'hfe00;
			16'hcc08: y = 16'hfe00;
			16'hcc09: y = 16'hfe00;
			16'hcc0a: y = 16'hfe00;
			16'hcc0b: y = 16'hfe00;
			16'hcc0c: y = 16'hfe00;
			16'hcc0d: y = 16'hfe00;
			16'hcc0e: y = 16'hfe00;
			16'hcc0f: y = 16'hfe00;
			16'hcc10: y = 16'hfe00;
			16'hcc11: y = 16'hfe00;
			16'hcc12: y = 16'hfe00;
			16'hcc13: y = 16'hfe00;
			16'hcc14: y = 16'hfe00;
			16'hcc15: y = 16'hfe00;
			16'hcc16: y = 16'hfe00;
			16'hcc17: y = 16'hfe00;
			16'hcc18: y = 16'hfe00;
			16'hcc19: y = 16'hfe00;
			16'hcc1a: y = 16'hfe00;
			16'hcc1b: y = 16'hfe00;
			16'hcc1c: y = 16'hfe00;
			16'hcc1d: y = 16'hfe00;
			16'hcc1e: y = 16'hfe00;
			16'hcc1f: y = 16'hfe00;
			16'hcc20: y = 16'hfe00;
			16'hcc21: y = 16'hfe00;
			16'hcc22: y = 16'hfe00;
			16'hcc23: y = 16'hfe00;
			16'hcc24: y = 16'hfe00;
			16'hcc25: y = 16'hfe00;
			16'hcc26: y = 16'hfe00;
			16'hcc27: y = 16'hfe00;
			16'hcc28: y = 16'hfe00;
			16'hcc29: y = 16'hfe00;
			16'hcc2a: y = 16'hfe00;
			16'hcc2b: y = 16'hfe00;
			16'hcc2c: y = 16'hfe00;
			16'hcc2d: y = 16'hfe00;
			16'hcc2e: y = 16'hfe00;
			16'hcc2f: y = 16'hfe00;
			16'hcc30: y = 16'hfe00;
			16'hcc31: y = 16'hfe00;
			16'hcc32: y = 16'hfe00;
			16'hcc33: y = 16'hfe00;
			16'hcc34: y = 16'hfe00;
			16'hcc35: y = 16'hfe00;
			16'hcc36: y = 16'hfe00;
			16'hcc37: y = 16'hfe00;
			16'hcc38: y = 16'hfe00;
			16'hcc39: y = 16'hfe00;
			16'hcc3a: y = 16'hfe00;
			16'hcc3b: y = 16'hfe00;
			16'hcc3c: y = 16'hfe00;
			16'hcc3d: y = 16'hfe00;
			16'hcc3e: y = 16'hfe00;
			16'hcc3f: y = 16'hfe00;
			16'hcc40: y = 16'hfe00;
			16'hcc41: y = 16'hfe00;
			16'hcc42: y = 16'hfe00;
			16'hcc43: y = 16'hfe00;
			16'hcc44: y = 16'hfe00;
			16'hcc45: y = 16'hfe00;
			16'hcc46: y = 16'hfe00;
			16'hcc47: y = 16'hfe00;
			16'hcc48: y = 16'hfe00;
			16'hcc49: y = 16'hfe00;
			16'hcc4a: y = 16'hfe00;
			16'hcc4b: y = 16'hfe00;
			16'hcc4c: y = 16'hfe00;
			16'hcc4d: y = 16'hfe00;
			16'hcc4e: y = 16'hfe00;
			16'hcc4f: y = 16'hfe00;
			16'hcc50: y = 16'hfe00;
			16'hcc51: y = 16'hfe00;
			16'hcc52: y = 16'hfe00;
			16'hcc53: y = 16'hfe00;
			16'hcc54: y = 16'hfe00;
			16'hcc55: y = 16'hfe00;
			16'hcc56: y = 16'hfe00;
			16'hcc57: y = 16'hfe00;
			16'hcc58: y = 16'hfe00;
			16'hcc59: y = 16'hfe00;
			16'hcc5a: y = 16'hfe00;
			16'hcc5b: y = 16'hfe00;
			16'hcc5c: y = 16'hfe00;
			16'hcc5d: y = 16'hfe00;
			16'hcc5e: y = 16'hfe00;
			16'hcc5f: y = 16'hfe00;
			16'hcc60: y = 16'hfe00;
			16'hcc61: y = 16'hfe00;
			16'hcc62: y = 16'hfe00;
			16'hcc63: y = 16'hfe00;
			16'hcc64: y = 16'hfe00;
			16'hcc65: y = 16'hfe00;
			16'hcc66: y = 16'hfe00;
			16'hcc67: y = 16'hfe00;
			16'hcc68: y = 16'hfe00;
			16'hcc69: y = 16'hfe00;
			16'hcc6a: y = 16'hfe00;
			16'hcc6b: y = 16'hfe00;
			16'hcc6c: y = 16'hfe00;
			16'hcc6d: y = 16'hfe00;
			16'hcc6e: y = 16'hfe00;
			16'hcc6f: y = 16'hfe00;
			16'hcc70: y = 16'hfe00;
			16'hcc71: y = 16'hfe00;
			16'hcc72: y = 16'hfe00;
			16'hcc73: y = 16'hfe00;
			16'hcc74: y = 16'hfe00;
			16'hcc75: y = 16'hfe00;
			16'hcc76: y = 16'hfe00;
			16'hcc77: y = 16'hfe00;
			16'hcc78: y = 16'hfe00;
			16'hcc79: y = 16'hfe00;
			16'hcc7a: y = 16'hfe00;
			16'hcc7b: y = 16'hfe00;
			16'hcc7c: y = 16'hfe00;
			16'hcc7d: y = 16'hfe00;
			16'hcc7e: y = 16'hfe00;
			16'hcc7f: y = 16'hfe00;
			16'hcc80: y = 16'hfe00;
			16'hcc81: y = 16'hfe00;
			16'hcc82: y = 16'hfe00;
			16'hcc83: y = 16'hfe00;
			16'hcc84: y = 16'hfe00;
			16'hcc85: y = 16'hfe00;
			16'hcc86: y = 16'hfe00;
			16'hcc87: y = 16'hfe00;
			16'hcc88: y = 16'hfe00;
			16'hcc89: y = 16'hfe00;
			16'hcc8a: y = 16'hfe00;
			16'hcc8b: y = 16'hfe00;
			16'hcc8c: y = 16'hfe00;
			16'hcc8d: y = 16'hfe00;
			16'hcc8e: y = 16'hfe00;
			16'hcc8f: y = 16'hfe00;
			16'hcc90: y = 16'hfe00;
			16'hcc91: y = 16'hfe00;
			16'hcc92: y = 16'hfe00;
			16'hcc93: y = 16'hfe00;
			16'hcc94: y = 16'hfe00;
			16'hcc95: y = 16'hfe00;
			16'hcc96: y = 16'hfe00;
			16'hcc97: y = 16'hfe00;
			16'hcc98: y = 16'hfe00;
			16'hcc99: y = 16'hfe00;
			16'hcc9a: y = 16'hfe00;
			16'hcc9b: y = 16'hfe00;
			16'hcc9c: y = 16'hfe00;
			16'hcc9d: y = 16'hfe00;
			16'hcc9e: y = 16'hfe00;
			16'hcc9f: y = 16'hfe00;
			16'hcca0: y = 16'hfe00;
			16'hcca1: y = 16'hfe00;
			16'hcca2: y = 16'hfe00;
			16'hcca3: y = 16'hfe00;
			16'hcca4: y = 16'hfe00;
			16'hcca5: y = 16'hfe00;
			16'hcca6: y = 16'hfe00;
			16'hcca7: y = 16'hfe00;
			16'hcca8: y = 16'hfe00;
			16'hcca9: y = 16'hfe00;
			16'hccaa: y = 16'hfe00;
			16'hccab: y = 16'hfe00;
			16'hccac: y = 16'hfe00;
			16'hccad: y = 16'hfe00;
			16'hccae: y = 16'hfe00;
			16'hccaf: y = 16'hfe00;
			16'hccb0: y = 16'hfe00;
			16'hccb1: y = 16'hfe00;
			16'hccb2: y = 16'hfe00;
			16'hccb3: y = 16'hfe00;
			16'hccb4: y = 16'hfe00;
			16'hccb5: y = 16'hfe00;
			16'hccb6: y = 16'hfe00;
			16'hccb7: y = 16'hfe00;
			16'hccb8: y = 16'hfe00;
			16'hccb9: y = 16'hfe00;
			16'hccba: y = 16'hfe00;
			16'hccbb: y = 16'hfe00;
			16'hccbc: y = 16'hfe00;
			16'hccbd: y = 16'hfe00;
			16'hccbe: y = 16'hfe00;
			16'hccbf: y = 16'hfe00;
			16'hccc0: y = 16'hfe00;
			16'hccc1: y = 16'hfe00;
			16'hccc2: y = 16'hfe00;
			16'hccc3: y = 16'hfe00;
			16'hccc4: y = 16'hfe00;
			16'hccc5: y = 16'hfe00;
			16'hccc6: y = 16'hfe00;
			16'hccc7: y = 16'hfe00;
			16'hccc8: y = 16'hfe00;
			16'hccc9: y = 16'hfe00;
			16'hccca: y = 16'hfe00;
			16'hcccb: y = 16'hfe00;
			16'hcccc: y = 16'hfe00;
			16'hcccd: y = 16'hfe00;
			16'hccce: y = 16'hfe00;
			16'hcccf: y = 16'hfe00;
			16'hccd0: y = 16'hfe00;
			16'hccd1: y = 16'hfe00;
			16'hccd2: y = 16'hfe00;
			16'hccd3: y = 16'hfe00;
			16'hccd4: y = 16'hfe00;
			16'hccd5: y = 16'hfe00;
			16'hccd6: y = 16'hfe00;
			16'hccd7: y = 16'hfe00;
			16'hccd8: y = 16'hfe00;
			16'hccd9: y = 16'hfe00;
			16'hccda: y = 16'hfe00;
			16'hccdb: y = 16'hfe00;
			16'hccdc: y = 16'hfe00;
			16'hccdd: y = 16'hfe00;
			16'hccde: y = 16'hfe00;
			16'hccdf: y = 16'hfe00;
			16'hcce0: y = 16'hfe00;
			16'hcce1: y = 16'hfe00;
			16'hcce2: y = 16'hfe00;
			16'hcce3: y = 16'hfe00;
			16'hcce4: y = 16'hfe00;
			16'hcce5: y = 16'hfe00;
			16'hcce6: y = 16'hfe00;
			16'hcce7: y = 16'hfe00;
			16'hcce8: y = 16'hfe00;
			16'hcce9: y = 16'hfe00;
			16'hccea: y = 16'hfe00;
			16'hcceb: y = 16'hfe00;
			16'hccec: y = 16'hfe00;
			16'hcced: y = 16'hfe00;
			16'hccee: y = 16'hfe00;
			16'hccef: y = 16'hfe00;
			16'hccf0: y = 16'hfe00;
			16'hccf1: y = 16'hfe00;
			16'hccf2: y = 16'hfe00;
			16'hccf3: y = 16'hfe00;
			16'hccf4: y = 16'hfe00;
			16'hccf5: y = 16'hfe00;
			16'hccf6: y = 16'hfe00;
			16'hccf7: y = 16'hfe00;
			16'hccf8: y = 16'hfe00;
			16'hccf9: y = 16'hfe00;
			16'hccfa: y = 16'hfe00;
			16'hccfb: y = 16'hfe00;
			16'hccfc: y = 16'hfe00;
			16'hccfd: y = 16'hfe00;
			16'hccfe: y = 16'hfe00;
			16'hccff: y = 16'hfe00;
			16'hcd00: y = 16'hfe00;
			16'hcd01: y = 16'hfe00;
			16'hcd02: y = 16'hfe00;
			16'hcd03: y = 16'hfe00;
			16'hcd04: y = 16'hfe00;
			16'hcd05: y = 16'hfe00;
			16'hcd06: y = 16'hfe00;
			16'hcd07: y = 16'hfe00;
			16'hcd08: y = 16'hfe00;
			16'hcd09: y = 16'hfe00;
			16'hcd0a: y = 16'hfe00;
			16'hcd0b: y = 16'hfe00;
			16'hcd0c: y = 16'hfe00;
			16'hcd0d: y = 16'hfe00;
			16'hcd0e: y = 16'hfe00;
			16'hcd0f: y = 16'hfe00;
			16'hcd10: y = 16'hfe00;
			16'hcd11: y = 16'hfe00;
			16'hcd12: y = 16'hfe00;
			16'hcd13: y = 16'hfe00;
			16'hcd14: y = 16'hfe00;
			16'hcd15: y = 16'hfe00;
			16'hcd16: y = 16'hfe00;
			16'hcd17: y = 16'hfe00;
			16'hcd18: y = 16'hfe00;
			16'hcd19: y = 16'hfe00;
			16'hcd1a: y = 16'hfe00;
			16'hcd1b: y = 16'hfe00;
			16'hcd1c: y = 16'hfe00;
			16'hcd1d: y = 16'hfe00;
			16'hcd1e: y = 16'hfe00;
			16'hcd1f: y = 16'hfe00;
			16'hcd20: y = 16'hfe00;
			16'hcd21: y = 16'hfe00;
			16'hcd22: y = 16'hfe00;
			16'hcd23: y = 16'hfe00;
			16'hcd24: y = 16'hfe00;
			16'hcd25: y = 16'hfe00;
			16'hcd26: y = 16'hfe00;
			16'hcd27: y = 16'hfe00;
			16'hcd28: y = 16'hfe00;
			16'hcd29: y = 16'hfe00;
			16'hcd2a: y = 16'hfe00;
			16'hcd2b: y = 16'hfe00;
			16'hcd2c: y = 16'hfe00;
			16'hcd2d: y = 16'hfe00;
			16'hcd2e: y = 16'hfe00;
			16'hcd2f: y = 16'hfe00;
			16'hcd30: y = 16'hfe00;
			16'hcd31: y = 16'hfe00;
			16'hcd32: y = 16'hfe00;
			16'hcd33: y = 16'hfe00;
			16'hcd34: y = 16'hfe00;
			16'hcd35: y = 16'hfe00;
			16'hcd36: y = 16'hfe00;
			16'hcd37: y = 16'hfe00;
			16'hcd38: y = 16'hfe00;
			16'hcd39: y = 16'hfe00;
			16'hcd3a: y = 16'hfe00;
			16'hcd3b: y = 16'hfe00;
			16'hcd3c: y = 16'hfe00;
			16'hcd3d: y = 16'hfe00;
			16'hcd3e: y = 16'hfe00;
			16'hcd3f: y = 16'hfe00;
			16'hcd40: y = 16'hfe00;
			16'hcd41: y = 16'hfe00;
			16'hcd42: y = 16'hfe00;
			16'hcd43: y = 16'hfe00;
			16'hcd44: y = 16'hfe00;
			16'hcd45: y = 16'hfe00;
			16'hcd46: y = 16'hfe00;
			16'hcd47: y = 16'hfe00;
			16'hcd48: y = 16'hfe00;
			16'hcd49: y = 16'hfe00;
			16'hcd4a: y = 16'hfe00;
			16'hcd4b: y = 16'hfe00;
			16'hcd4c: y = 16'hfe00;
			16'hcd4d: y = 16'hfe00;
			16'hcd4e: y = 16'hfe00;
			16'hcd4f: y = 16'hfe00;
			16'hcd50: y = 16'hfe00;
			16'hcd51: y = 16'hfe00;
			16'hcd52: y = 16'hfe00;
			16'hcd53: y = 16'hfe00;
			16'hcd54: y = 16'hfe00;
			16'hcd55: y = 16'hfe00;
			16'hcd56: y = 16'hfe00;
			16'hcd57: y = 16'hfe00;
			16'hcd58: y = 16'hfe00;
			16'hcd59: y = 16'hfe00;
			16'hcd5a: y = 16'hfe00;
			16'hcd5b: y = 16'hfe00;
			16'hcd5c: y = 16'hfe00;
			16'hcd5d: y = 16'hfe00;
			16'hcd5e: y = 16'hfe00;
			16'hcd5f: y = 16'hfe00;
			16'hcd60: y = 16'hfe00;
			16'hcd61: y = 16'hfe00;
			16'hcd62: y = 16'hfe00;
			16'hcd63: y = 16'hfe00;
			16'hcd64: y = 16'hfe00;
			16'hcd65: y = 16'hfe00;
			16'hcd66: y = 16'hfe00;
			16'hcd67: y = 16'hfe00;
			16'hcd68: y = 16'hfe00;
			16'hcd69: y = 16'hfe00;
			16'hcd6a: y = 16'hfe00;
			16'hcd6b: y = 16'hfe00;
			16'hcd6c: y = 16'hfe00;
			16'hcd6d: y = 16'hfe00;
			16'hcd6e: y = 16'hfe00;
			16'hcd6f: y = 16'hfe00;
			16'hcd70: y = 16'hfe00;
			16'hcd71: y = 16'hfe00;
			16'hcd72: y = 16'hfe00;
			16'hcd73: y = 16'hfe00;
			16'hcd74: y = 16'hfe00;
			16'hcd75: y = 16'hfe00;
			16'hcd76: y = 16'hfe00;
			16'hcd77: y = 16'hfe00;
			16'hcd78: y = 16'hfe00;
			16'hcd79: y = 16'hfe00;
			16'hcd7a: y = 16'hfe00;
			16'hcd7b: y = 16'hfe00;
			16'hcd7c: y = 16'hfe00;
			16'hcd7d: y = 16'hfe00;
			16'hcd7e: y = 16'hfe00;
			16'hcd7f: y = 16'hfe00;
			16'hcd80: y = 16'hfe00;
			16'hcd81: y = 16'hfe00;
			16'hcd82: y = 16'hfe00;
			16'hcd83: y = 16'hfe00;
			16'hcd84: y = 16'hfe00;
			16'hcd85: y = 16'hfe00;
			16'hcd86: y = 16'hfe00;
			16'hcd87: y = 16'hfe00;
			16'hcd88: y = 16'hfe00;
			16'hcd89: y = 16'hfe00;
			16'hcd8a: y = 16'hfe00;
			16'hcd8b: y = 16'hfe00;
			16'hcd8c: y = 16'hfe00;
			16'hcd8d: y = 16'hfe00;
			16'hcd8e: y = 16'hfe00;
			16'hcd8f: y = 16'hfe00;
			16'hcd90: y = 16'hfe00;
			16'hcd91: y = 16'hfe00;
			16'hcd92: y = 16'hfe00;
			16'hcd93: y = 16'hfe00;
			16'hcd94: y = 16'hfe00;
			16'hcd95: y = 16'hfe00;
			16'hcd96: y = 16'hfe00;
			16'hcd97: y = 16'hfe00;
			16'hcd98: y = 16'hfe00;
			16'hcd99: y = 16'hfe00;
			16'hcd9a: y = 16'hfe00;
			16'hcd9b: y = 16'hfe00;
			16'hcd9c: y = 16'hfe00;
			16'hcd9d: y = 16'hfe00;
			16'hcd9e: y = 16'hfe00;
			16'hcd9f: y = 16'hfe00;
			16'hcda0: y = 16'hfe00;
			16'hcda1: y = 16'hfe00;
			16'hcda2: y = 16'hfe00;
			16'hcda3: y = 16'hfe00;
			16'hcda4: y = 16'hfe00;
			16'hcda5: y = 16'hfe00;
			16'hcda6: y = 16'hfe00;
			16'hcda7: y = 16'hfe00;
			16'hcda8: y = 16'hfe00;
			16'hcda9: y = 16'hfe00;
			16'hcdaa: y = 16'hfe00;
			16'hcdab: y = 16'hfe00;
			16'hcdac: y = 16'hfe00;
			16'hcdad: y = 16'hfe00;
			16'hcdae: y = 16'hfe00;
			16'hcdaf: y = 16'hfe00;
			16'hcdb0: y = 16'hfe00;
			16'hcdb1: y = 16'hfe00;
			16'hcdb2: y = 16'hfe00;
			16'hcdb3: y = 16'hfe00;
			16'hcdb4: y = 16'hfe00;
			16'hcdb5: y = 16'hfe00;
			16'hcdb6: y = 16'hfe00;
			16'hcdb7: y = 16'hfe00;
			16'hcdb8: y = 16'hfe00;
			16'hcdb9: y = 16'hfe00;
			16'hcdba: y = 16'hfe00;
			16'hcdbb: y = 16'hfe00;
			16'hcdbc: y = 16'hfe00;
			16'hcdbd: y = 16'hfe00;
			16'hcdbe: y = 16'hfe00;
			16'hcdbf: y = 16'hfe00;
			16'hcdc0: y = 16'hfe00;
			16'hcdc1: y = 16'hfe00;
			16'hcdc2: y = 16'hfe00;
			16'hcdc3: y = 16'hfe00;
			16'hcdc4: y = 16'hfe00;
			16'hcdc5: y = 16'hfe00;
			16'hcdc6: y = 16'hfe00;
			16'hcdc7: y = 16'hfe00;
			16'hcdc8: y = 16'hfe00;
			16'hcdc9: y = 16'hfe00;
			16'hcdca: y = 16'hfe00;
			16'hcdcb: y = 16'hfe00;
			16'hcdcc: y = 16'hfe00;
			16'hcdcd: y = 16'hfe00;
			16'hcdce: y = 16'hfe00;
			16'hcdcf: y = 16'hfe00;
			16'hcdd0: y = 16'hfe00;
			16'hcdd1: y = 16'hfe00;
			16'hcdd2: y = 16'hfe00;
			16'hcdd3: y = 16'hfe00;
			16'hcdd4: y = 16'hfe00;
			16'hcdd5: y = 16'hfe00;
			16'hcdd6: y = 16'hfe00;
			16'hcdd7: y = 16'hfe00;
			16'hcdd8: y = 16'hfe00;
			16'hcdd9: y = 16'hfe00;
			16'hcdda: y = 16'hfe00;
			16'hcddb: y = 16'hfe00;
			16'hcddc: y = 16'hfe00;
			16'hcddd: y = 16'hfe00;
			16'hcdde: y = 16'hfe00;
			16'hcddf: y = 16'hfe00;
			16'hcde0: y = 16'hfe00;
			16'hcde1: y = 16'hfe00;
			16'hcde2: y = 16'hfe00;
			16'hcde3: y = 16'hfe00;
			16'hcde4: y = 16'hfe00;
			16'hcde5: y = 16'hfe00;
			16'hcde6: y = 16'hfe00;
			16'hcde7: y = 16'hfe00;
			16'hcde8: y = 16'hfe00;
			16'hcde9: y = 16'hfe00;
			16'hcdea: y = 16'hfe00;
			16'hcdeb: y = 16'hfe00;
			16'hcdec: y = 16'hfe00;
			16'hcded: y = 16'hfe00;
			16'hcdee: y = 16'hfe00;
			16'hcdef: y = 16'hfe00;
			16'hcdf0: y = 16'hfe00;
			16'hcdf1: y = 16'hfe00;
			16'hcdf2: y = 16'hfe00;
			16'hcdf3: y = 16'hfe00;
			16'hcdf4: y = 16'hfe00;
			16'hcdf5: y = 16'hfe00;
			16'hcdf6: y = 16'hfe00;
			16'hcdf7: y = 16'hfe00;
			16'hcdf8: y = 16'hfe00;
			16'hcdf9: y = 16'hfe00;
			16'hcdfa: y = 16'hfe00;
			16'hcdfb: y = 16'hfe00;
			16'hcdfc: y = 16'hfe00;
			16'hcdfd: y = 16'hfe00;
			16'hcdfe: y = 16'hfe00;
			16'hcdff: y = 16'hfe00;
			16'hce00: y = 16'hfe00;
			16'hce01: y = 16'hfe00;
			16'hce02: y = 16'hfe00;
			16'hce03: y = 16'hfe00;
			16'hce04: y = 16'hfe00;
			16'hce05: y = 16'hfe00;
			16'hce06: y = 16'hfe00;
			16'hce07: y = 16'hfe00;
			16'hce08: y = 16'hfe00;
			16'hce09: y = 16'hfe00;
			16'hce0a: y = 16'hfe00;
			16'hce0b: y = 16'hfe00;
			16'hce0c: y = 16'hfe00;
			16'hce0d: y = 16'hfe00;
			16'hce0e: y = 16'hfe00;
			16'hce0f: y = 16'hfe00;
			16'hce10: y = 16'hfe00;
			16'hce11: y = 16'hfe00;
			16'hce12: y = 16'hfe00;
			16'hce13: y = 16'hfe00;
			16'hce14: y = 16'hfe00;
			16'hce15: y = 16'hfe00;
			16'hce16: y = 16'hfe00;
			16'hce17: y = 16'hfe00;
			16'hce18: y = 16'hfe00;
			16'hce19: y = 16'hfe00;
			16'hce1a: y = 16'hfe00;
			16'hce1b: y = 16'hfe00;
			16'hce1c: y = 16'hfe00;
			16'hce1d: y = 16'hfe00;
			16'hce1e: y = 16'hfe00;
			16'hce1f: y = 16'hfe00;
			16'hce20: y = 16'hfe00;
			16'hce21: y = 16'hfe00;
			16'hce22: y = 16'hfe00;
			16'hce23: y = 16'hfe00;
			16'hce24: y = 16'hfe00;
			16'hce25: y = 16'hfe00;
			16'hce26: y = 16'hfe00;
			16'hce27: y = 16'hfe00;
			16'hce28: y = 16'hfe00;
			16'hce29: y = 16'hfe00;
			16'hce2a: y = 16'hfe00;
			16'hce2b: y = 16'hfe00;
			16'hce2c: y = 16'hfe00;
			16'hce2d: y = 16'hfe00;
			16'hce2e: y = 16'hfe00;
			16'hce2f: y = 16'hfe00;
			16'hce30: y = 16'hfe00;
			16'hce31: y = 16'hfe00;
			16'hce32: y = 16'hfe00;
			16'hce33: y = 16'hfe00;
			16'hce34: y = 16'hfe00;
			16'hce35: y = 16'hfe00;
			16'hce36: y = 16'hfe00;
			16'hce37: y = 16'hfe00;
			16'hce38: y = 16'hfe00;
			16'hce39: y = 16'hfe00;
			16'hce3a: y = 16'hfe00;
			16'hce3b: y = 16'hfe00;
			16'hce3c: y = 16'hfe00;
			16'hce3d: y = 16'hfe00;
			16'hce3e: y = 16'hfe00;
			16'hce3f: y = 16'hfe00;
			16'hce40: y = 16'hfe00;
			16'hce41: y = 16'hfe00;
			16'hce42: y = 16'hfe00;
			16'hce43: y = 16'hfe00;
			16'hce44: y = 16'hfe00;
			16'hce45: y = 16'hfe00;
			16'hce46: y = 16'hfe00;
			16'hce47: y = 16'hfe00;
			16'hce48: y = 16'hfe00;
			16'hce49: y = 16'hfe00;
			16'hce4a: y = 16'hfe00;
			16'hce4b: y = 16'hfe00;
			16'hce4c: y = 16'hfe00;
			16'hce4d: y = 16'hfe00;
			16'hce4e: y = 16'hfe00;
			16'hce4f: y = 16'hfe00;
			16'hce50: y = 16'hfe00;
			16'hce51: y = 16'hfe00;
			16'hce52: y = 16'hfe00;
			16'hce53: y = 16'hfe00;
			16'hce54: y = 16'hfe00;
			16'hce55: y = 16'hfe00;
			16'hce56: y = 16'hfe00;
			16'hce57: y = 16'hfe00;
			16'hce58: y = 16'hfe00;
			16'hce59: y = 16'hfe00;
			16'hce5a: y = 16'hfe00;
			16'hce5b: y = 16'hfe00;
			16'hce5c: y = 16'hfe00;
			16'hce5d: y = 16'hfe00;
			16'hce5e: y = 16'hfe00;
			16'hce5f: y = 16'hfe00;
			16'hce60: y = 16'hfe00;
			16'hce61: y = 16'hfe00;
			16'hce62: y = 16'hfe00;
			16'hce63: y = 16'hfe00;
			16'hce64: y = 16'hfe00;
			16'hce65: y = 16'hfe00;
			16'hce66: y = 16'hfe00;
			16'hce67: y = 16'hfe00;
			16'hce68: y = 16'hfe00;
			16'hce69: y = 16'hfe00;
			16'hce6a: y = 16'hfe00;
			16'hce6b: y = 16'hfe00;
			16'hce6c: y = 16'hfe00;
			16'hce6d: y = 16'hfe00;
			16'hce6e: y = 16'hfe00;
			16'hce6f: y = 16'hfe00;
			16'hce70: y = 16'hfe00;
			16'hce71: y = 16'hfe00;
			16'hce72: y = 16'hfe00;
			16'hce73: y = 16'hfe00;
			16'hce74: y = 16'hfe00;
			16'hce75: y = 16'hfe00;
			16'hce76: y = 16'hfe00;
			16'hce77: y = 16'hfe00;
			16'hce78: y = 16'hfe00;
			16'hce79: y = 16'hfe00;
			16'hce7a: y = 16'hfe00;
			16'hce7b: y = 16'hfe00;
			16'hce7c: y = 16'hfe00;
			16'hce7d: y = 16'hfe00;
			16'hce7e: y = 16'hfe00;
			16'hce7f: y = 16'hfe00;
			16'hce80: y = 16'hfe00;
			16'hce81: y = 16'hfe00;
			16'hce82: y = 16'hfe00;
			16'hce83: y = 16'hfe00;
			16'hce84: y = 16'hfe00;
			16'hce85: y = 16'hfe00;
			16'hce86: y = 16'hfe00;
			16'hce87: y = 16'hfe00;
			16'hce88: y = 16'hfe00;
			16'hce89: y = 16'hfe00;
			16'hce8a: y = 16'hfe00;
			16'hce8b: y = 16'hfe00;
			16'hce8c: y = 16'hfe00;
			16'hce8d: y = 16'hfe00;
			16'hce8e: y = 16'hfe00;
			16'hce8f: y = 16'hfe00;
			16'hce90: y = 16'hfe00;
			16'hce91: y = 16'hfe00;
			16'hce92: y = 16'hfe00;
			16'hce93: y = 16'hfe00;
			16'hce94: y = 16'hfe00;
			16'hce95: y = 16'hfe00;
			16'hce96: y = 16'hfe00;
			16'hce97: y = 16'hfe00;
			16'hce98: y = 16'hfe00;
			16'hce99: y = 16'hfe00;
			16'hce9a: y = 16'hfe00;
			16'hce9b: y = 16'hfe00;
			16'hce9c: y = 16'hfe00;
			16'hce9d: y = 16'hfe00;
			16'hce9e: y = 16'hfe00;
			16'hce9f: y = 16'hfe00;
			16'hcea0: y = 16'hfe00;
			16'hcea1: y = 16'hfe00;
			16'hcea2: y = 16'hfe00;
			16'hcea3: y = 16'hfe00;
			16'hcea4: y = 16'hfe00;
			16'hcea5: y = 16'hfe00;
			16'hcea6: y = 16'hfe00;
			16'hcea7: y = 16'hfe00;
			16'hcea8: y = 16'hfe00;
			16'hcea9: y = 16'hfe00;
			16'hceaa: y = 16'hfe00;
			16'hceab: y = 16'hfe00;
			16'hceac: y = 16'hfe00;
			16'hcead: y = 16'hfe00;
			16'hceae: y = 16'hfe00;
			16'hceaf: y = 16'hfe00;
			16'hceb0: y = 16'hfe00;
			16'hceb1: y = 16'hfe00;
			16'hceb2: y = 16'hfe00;
			16'hceb3: y = 16'hfe00;
			16'hceb4: y = 16'hfe00;
			16'hceb5: y = 16'hfe00;
			16'hceb6: y = 16'hfe00;
			16'hceb7: y = 16'hfe00;
			16'hceb8: y = 16'hfe00;
			16'hceb9: y = 16'hfe00;
			16'hceba: y = 16'hfe00;
			16'hcebb: y = 16'hfe00;
			16'hcebc: y = 16'hfe00;
			16'hcebd: y = 16'hfe00;
			16'hcebe: y = 16'hfe00;
			16'hcebf: y = 16'hfe00;
			16'hcec0: y = 16'hfe00;
			16'hcec1: y = 16'hfe00;
			16'hcec2: y = 16'hfe00;
			16'hcec3: y = 16'hfe00;
			16'hcec4: y = 16'hfe00;
			16'hcec5: y = 16'hfe00;
			16'hcec6: y = 16'hfe00;
			16'hcec7: y = 16'hfe00;
			16'hcec8: y = 16'hfe00;
			16'hcec9: y = 16'hfe00;
			16'hceca: y = 16'hfe00;
			16'hcecb: y = 16'hfe00;
			16'hcecc: y = 16'hfe00;
			16'hcecd: y = 16'hfe00;
			16'hcece: y = 16'hfe00;
			16'hcecf: y = 16'hfe00;
			16'hced0: y = 16'hfe00;
			16'hced1: y = 16'hfe00;
			16'hced2: y = 16'hfe00;
			16'hced3: y = 16'hfe00;
			16'hced4: y = 16'hfe00;
			16'hced5: y = 16'hfe00;
			16'hced6: y = 16'hfe00;
			16'hced7: y = 16'hfe00;
			16'hced8: y = 16'hfe00;
			16'hced9: y = 16'hfe00;
			16'hceda: y = 16'hfe00;
			16'hcedb: y = 16'hfe00;
			16'hcedc: y = 16'hfe00;
			16'hcedd: y = 16'hfe00;
			16'hcede: y = 16'hfe00;
			16'hcedf: y = 16'hfe00;
			16'hcee0: y = 16'hfe00;
			16'hcee1: y = 16'hfe00;
			16'hcee2: y = 16'hfe00;
			16'hcee3: y = 16'hfe00;
			16'hcee4: y = 16'hfe00;
			16'hcee5: y = 16'hfe00;
			16'hcee6: y = 16'hfe00;
			16'hcee7: y = 16'hfe00;
			16'hcee8: y = 16'hfe00;
			16'hcee9: y = 16'hfe00;
			16'hceea: y = 16'hfe00;
			16'hceeb: y = 16'hfe00;
			16'hceec: y = 16'hfe00;
			16'hceed: y = 16'hfe00;
			16'hceee: y = 16'hfe00;
			16'hceef: y = 16'hfe00;
			16'hcef0: y = 16'hfe00;
			16'hcef1: y = 16'hfe00;
			16'hcef2: y = 16'hfe00;
			16'hcef3: y = 16'hfe00;
			16'hcef4: y = 16'hfe00;
			16'hcef5: y = 16'hfe00;
			16'hcef6: y = 16'hfe00;
			16'hcef7: y = 16'hfe00;
			16'hcef8: y = 16'hfe00;
			16'hcef9: y = 16'hfe00;
			16'hcefa: y = 16'hfe00;
			16'hcefb: y = 16'hfe00;
			16'hcefc: y = 16'hfe00;
			16'hcefd: y = 16'hfe00;
			16'hcefe: y = 16'hfe00;
			16'hceff: y = 16'hfe00;
			16'hcf00: y = 16'hfe00;
			16'hcf01: y = 16'hfe00;
			16'hcf02: y = 16'hfe00;
			16'hcf03: y = 16'hfe00;
			16'hcf04: y = 16'hfe00;
			16'hcf05: y = 16'hfe00;
			16'hcf06: y = 16'hfe00;
			16'hcf07: y = 16'hfe00;
			16'hcf08: y = 16'hfe00;
			16'hcf09: y = 16'hfe00;
			16'hcf0a: y = 16'hfe00;
			16'hcf0b: y = 16'hfe00;
			16'hcf0c: y = 16'hfe00;
			16'hcf0d: y = 16'hfe00;
			16'hcf0e: y = 16'hfe00;
			16'hcf0f: y = 16'hfe00;
			16'hcf10: y = 16'hfe00;
			16'hcf11: y = 16'hfe00;
			16'hcf12: y = 16'hfe00;
			16'hcf13: y = 16'hfe00;
			16'hcf14: y = 16'hfe00;
			16'hcf15: y = 16'hfe00;
			16'hcf16: y = 16'hfe00;
			16'hcf17: y = 16'hfe00;
			16'hcf18: y = 16'hfe00;
			16'hcf19: y = 16'hfe00;
			16'hcf1a: y = 16'hfe00;
			16'hcf1b: y = 16'hfe00;
			16'hcf1c: y = 16'hfe00;
			16'hcf1d: y = 16'hfe00;
			16'hcf1e: y = 16'hfe00;
			16'hcf1f: y = 16'hfe00;
			16'hcf20: y = 16'hfe00;
			16'hcf21: y = 16'hfe00;
			16'hcf22: y = 16'hfe00;
			16'hcf23: y = 16'hfe00;
			16'hcf24: y = 16'hfe00;
			16'hcf25: y = 16'hfe00;
			16'hcf26: y = 16'hfe00;
			16'hcf27: y = 16'hfe00;
			16'hcf28: y = 16'hfe00;
			16'hcf29: y = 16'hfe00;
			16'hcf2a: y = 16'hfe00;
			16'hcf2b: y = 16'hfe00;
			16'hcf2c: y = 16'hfe00;
			16'hcf2d: y = 16'hfe00;
			16'hcf2e: y = 16'hfe00;
			16'hcf2f: y = 16'hfe00;
			16'hcf30: y = 16'hfe00;
			16'hcf31: y = 16'hfe00;
			16'hcf32: y = 16'hfe00;
			16'hcf33: y = 16'hfe00;
			16'hcf34: y = 16'hfe00;
			16'hcf35: y = 16'hfe00;
			16'hcf36: y = 16'hfe00;
			16'hcf37: y = 16'hfe00;
			16'hcf38: y = 16'hfe00;
			16'hcf39: y = 16'hfe00;
			16'hcf3a: y = 16'hfe00;
			16'hcf3b: y = 16'hfe00;
			16'hcf3c: y = 16'hfe00;
			16'hcf3d: y = 16'hfe00;
			16'hcf3e: y = 16'hfe00;
			16'hcf3f: y = 16'hfe00;
			16'hcf40: y = 16'hfe00;
			16'hcf41: y = 16'hfe00;
			16'hcf42: y = 16'hfe00;
			16'hcf43: y = 16'hfe00;
			16'hcf44: y = 16'hfe00;
			16'hcf45: y = 16'hfe00;
			16'hcf46: y = 16'hfe00;
			16'hcf47: y = 16'hfe00;
			16'hcf48: y = 16'hfe00;
			16'hcf49: y = 16'hfe00;
			16'hcf4a: y = 16'hfe00;
			16'hcf4b: y = 16'hfe00;
			16'hcf4c: y = 16'hfe00;
			16'hcf4d: y = 16'hfe00;
			16'hcf4e: y = 16'hfe00;
			16'hcf4f: y = 16'hfe00;
			16'hcf50: y = 16'hfe00;
			16'hcf51: y = 16'hfe00;
			16'hcf52: y = 16'hfe00;
			16'hcf53: y = 16'hfe00;
			16'hcf54: y = 16'hfe00;
			16'hcf55: y = 16'hfe00;
			16'hcf56: y = 16'hfe00;
			16'hcf57: y = 16'hfe00;
			16'hcf58: y = 16'hfe00;
			16'hcf59: y = 16'hfe00;
			16'hcf5a: y = 16'hfe00;
			16'hcf5b: y = 16'hfe00;
			16'hcf5c: y = 16'hfe00;
			16'hcf5d: y = 16'hfe00;
			16'hcf5e: y = 16'hfe00;
			16'hcf5f: y = 16'hfe00;
			16'hcf60: y = 16'hfe00;
			16'hcf61: y = 16'hfe00;
			16'hcf62: y = 16'hfe00;
			16'hcf63: y = 16'hfe00;
			16'hcf64: y = 16'hfe00;
			16'hcf65: y = 16'hfe00;
			16'hcf66: y = 16'hfe00;
			16'hcf67: y = 16'hfe00;
			16'hcf68: y = 16'hfe00;
			16'hcf69: y = 16'hfe00;
			16'hcf6a: y = 16'hfe00;
			16'hcf6b: y = 16'hfe00;
			16'hcf6c: y = 16'hfe00;
			16'hcf6d: y = 16'hfe00;
			16'hcf6e: y = 16'hfe00;
			16'hcf6f: y = 16'hfe00;
			16'hcf70: y = 16'hfe00;
			16'hcf71: y = 16'hfe00;
			16'hcf72: y = 16'hfe00;
			16'hcf73: y = 16'hfe00;
			16'hcf74: y = 16'hfe00;
			16'hcf75: y = 16'hfe00;
			16'hcf76: y = 16'hfe00;
			16'hcf77: y = 16'hfe00;
			16'hcf78: y = 16'hfe00;
			16'hcf79: y = 16'hfe00;
			16'hcf7a: y = 16'hfe00;
			16'hcf7b: y = 16'hfe00;
			16'hcf7c: y = 16'hfe00;
			16'hcf7d: y = 16'hfe00;
			16'hcf7e: y = 16'hfe00;
			16'hcf7f: y = 16'hfe00;
			16'hcf80: y = 16'hfe00;
			16'hcf81: y = 16'hfe00;
			16'hcf82: y = 16'hfe00;
			16'hcf83: y = 16'hfe00;
			16'hcf84: y = 16'hfe00;
			16'hcf85: y = 16'hfe00;
			16'hcf86: y = 16'hfe00;
			16'hcf87: y = 16'hfe00;
			16'hcf88: y = 16'hfe00;
			16'hcf89: y = 16'hfe00;
			16'hcf8a: y = 16'hfe00;
			16'hcf8b: y = 16'hfe00;
			16'hcf8c: y = 16'hfe00;
			16'hcf8d: y = 16'hfe00;
			16'hcf8e: y = 16'hfe00;
			16'hcf8f: y = 16'hfe00;
			16'hcf90: y = 16'hfe00;
			16'hcf91: y = 16'hfe00;
			16'hcf92: y = 16'hfe00;
			16'hcf93: y = 16'hfe00;
			16'hcf94: y = 16'hfe00;
			16'hcf95: y = 16'hfe00;
			16'hcf96: y = 16'hfe00;
			16'hcf97: y = 16'hfe00;
			16'hcf98: y = 16'hfe00;
			16'hcf99: y = 16'hfe00;
			16'hcf9a: y = 16'hfe00;
			16'hcf9b: y = 16'hfe00;
			16'hcf9c: y = 16'hfe00;
			16'hcf9d: y = 16'hfe00;
			16'hcf9e: y = 16'hfe00;
			16'hcf9f: y = 16'hfe00;
			16'hcfa0: y = 16'hfe00;
			16'hcfa1: y = 16'hfe00;
			16'hcfa2: y = 16'hfe00;
			16'hcfa3: y = 16'hfe00;
			16'hcfa4: y = 16'hfe00;
			16'hcfa5: y = 16'hfe00;
			16'hcfa6: y = 16'hfe00;
			16'hcfa7: y = 16'hfe00;
			16'hcfa8: y = 16'hfe00;
			16'hcfa9: y = 16'hfe00;
			16'hcfaa: y = 16'hfe00;
			16'hcfab: y = 16'hfe00;
			16'hcfac: y = 16'hfe00;
			16'hcfad: y = 16'hfe00;
			16'hcfae: y = 16'hfe00;
			16'hcfaf: y = 16'hfe00;
			16'hcfb0: y = 16'hfe00;
			16'hcfb1: y = 16'hfe00;
			16'hcfb2: y = 16'hfe00;
			16'hcfb3: y = 16'hfe00;
			16'hcfb4: y = 16'hfe00;
			16'hcfb5: y = 16'hfe00;
			16'hcfb6: y = 16'hfe00;
			16'hcfb7: y = 16'hfe00;
			16'hcfb8: y = 16'hfe00;
			16'hcfb9: y = 16'hfe00;
			16'hcfba: y = 16'hfe00;
			16'hcfbb: y = 16'hfe00;
			16'hcfbc: y = 16'hfe00;
			16'hcfbd: y = 16'hfe00;
			16'hcfbe: y = 16'hfe00;
			16'hcfbf: y = 16'hfe00;
			16'hcfc0: y = 16'hfe00;
			16'hcfc1: y = 16'hfe00;
			16'hcfc2: y = 16'hfe00;
			16'hcfc3: y = 16'hfe00;
			16'hcfc4: y = 16'hfe00;
			16'hcfc5: y = 16'hfe00;
			16'hcfc6: y = 16'hfe00;
			16'hcfc7: y = 16'hfe00;
			16'hcfc8: y = 16'hfe00;
			16'hcfc9: y = 16'hfe00;
			16'hcfca: y = 16'hfe00;
			16'hcfcb: y = 16'hfe00;
			16'hcfcc: y = 16'hfe00;
			16'hcfcd: y = 16'hfe00;
			16'hcfce: y = 16'hfe00;
			16'hcfcf: y = 16'hfe00;
			16'hcfd0: y = 16'hfe00;
			16'hcfd1: y = 16'hfe00;
			16'hcfd2: y = 16'hfe00;
			16'hcfd3: y = 16'hfe00;
			16'hcfd4: y = 16'hfe00;
			16'hcfd5: y = 16'hfe00;
			16'hcfd6: y = 16'hfe00;
			16'hcfd7: y = 16'hfe00;
			16'hcfd8: y = 16'hfe00;
			16'hcfd9: y = 16'hfe00;
			16'hcfda: y = 16'hfe00;
			16'hcfdb: y = 16'hfe00;
			16'hcfdc: y = 16'hfe00;
			16'hcfdd: y = 16'hfe00;
			16'hcfde: y = 16'hfe00;
			16'hcfdf: y = 16'hfe00;
			16'hcfe0: y = 16'hfe00;
			16'hcfe1: y = 16'hfe00;
			16'hcfe2: y = 16'hfe00;
			16'hcfe3: y = 16'hfe00;
			16'hcfe4: y = 16'hfe00;
			16'hcfe5: y = 16'hfe00;
			16'hcfe6: y = 16'hfe00;
			16'hcfe7: y = 16'hfe00;
			16'hcfe8: y = 16'hfe00;
			16'hcfe9: y = 16'hfe00;
			16'hcfea: y = 16'hfe00;
			16'hcfeb: y = 16'hfe00;
			16'hcfec: y = 16'hfe00;
			16'hcfed: y = 16'hfe00;
			16'hcfee: y = 16'hfe00;
			16'hcfef: y = 16'hfe00;
			16'hcff0: y = 16'hfe00;
			16'hcff1: y = 16'hfe00;
			16'hcff2: y = 16'hfe00;
			16'hcff3: y = 16'hfe00;
			16'hcff4: y = 16'hfe00;
			16'hcff5: y = 16'hfe00;
			16'hcff6: y = 16'hfe00;
			16'hcff7: y = 16'hfe00;
			16'hcff8: y = 16'hfe00;
			16'hcff9: y = 16'hfe00;
			16'hcffa: y = 16'hfe00;
			16'hcffb: y = 16'hfe00;
			16'hcffc: y = 16'hfe00;
			16'hcffd: y = 16'hfe00;
			16'hcffe: y = 16'hfe00;
			16'hcfff: y = 16'hfe00;
			16'hd000: y = 16'hfe00;
			16'hd001: y = 16'hfe00;
			16'hd002: y = 16'hfe00;
			16'hd003: y = 16'hfe00;
			16'hd004: y = 16'hfe00;
			16'hd005: y = 16'hfe00;
			16'hd006: y = 16'hfe00;
			16'hd007: y = 16'hfe00;
			16'hd008: y = 16'hfe00;
			16'hd009: y = 16'hfe00;
			16'hd00a: y = 16'hfe00;
			16'hd00b: y = 16'hfe00;
			16'hd00c: y = 16'hfe00;
			16'hd00d: y = 16'hfe00;
			16'hd00e: y = 16'hfe00;
			16'hd00f: y = 16'hfe00;
			16'hd010: y = 16'hfe00;
			16'hd011: y = 16'hfe00;
			16'hd012: y = 16'hfe00;
			16'hd013: y = 16'hfe00;
			16'hd014: y = 16'hfe00;
			16'hd015: y = 16'hfe00;
			16'hd016: y = 16'hfe00;
			16'hd017: y = 16'hfe00;
			16'hd018: y = 16'hfe00;
			16'hd019: y = 16'hfe00;
			16'hd01a: y = 16'hfe00;
			16'hd01b: y = 16'hfe00;
			16'hd01c: y = 16'hfe00;
			16'hd01d: y = 16'hfe00;
			16'hd01e: y = 16'hfe00;
			16'hd01f: y = 16'hfe00;
			16'hd020: y = 16'hfe00;
			16'hd021: y = 16'hfe00;
			16'hd022: y = 16'hfe00;
			16'hd023: y = 16'hfe00;
			16'hd024: y = 16'hfe00;
			16'hd025: y = 16'hfe00;
			16'hd026: y = 16'hfe00;
			16'hd027: y = 16'hfe00;
			16'hd028: y = 16'hfe00;
			16'hd029: y = 16'hfe00;
			16'hd02a: y = 16'hfe00;
			16'hd02b: y = 16'hfe00;
			16'hd02c: y = 16'hfe00;
			16'hd02d: y = 16'hfe00;
			16'hd02e: y = 16'hfe00;
			16'hd02f: y = 16'hfe00;
			16'hd030: y = 16'hfe00;
			16'hd031: y = 16'hfe00;
			16'hd032: y = 16'hfe00;
			16'hd033: y = 16'hfe00;
			16'hd034: y = 16'hfe00;
			16'hd035: y = 16'hfe00;
			16'hd036: y = 16'hfe00;
			16'hd037: y = 16'hfe00;
			16'hd038: y = 16'hfe00;
			16'hd039: y = 16'hfe00;
			16'hd03a: y = 16'hfe00;
			16'hd03b: y = 16'hfe00;
			16'hd03c: y = 16'hfe00;
			16'hd03d: y = 16'hfe00;
			16'hd03e: y = 16'hfe00;
			16'hd03f: y = 16'hfe00;
			16'hd040: y = 16'hfe00;
			16'hd041: y = 16'hfe00;
			16'hd042: y = 16'hfe00;
			16'hd043: y = 16'hfe00;
			16'hd044: y = 16'hfe00;
			16'hd045: y = 16'hfe00;
			16'hd046: y = 16'hfe00;
			16'hd047: y = 16'hfe00;
			16'hd048: y = 16'hfe00;
			16'hd049: y = 16'hfe00;
			16'hd04a: y = 16'hfe00;
			16'hd04b: y = 16'hfe00;
			16'hd04c: y = 16'hfe00;
			16'hd04d: y = 16'hfe00;
			16'hd04e: y = 16'hfe00;
			16'hd04f: y = 16'hfe00;
			16'hd050: y = 16'hfe00;
			16'hd051: y = 16'hfe00;
			16'hd052: y = 16'hfe00;
			16'hd053: y = 16'hfe00;
			16'hd054: y = 16'hfe00;
			16'hd055: y = 16'hfe00;
			16'hd056: y = 16'hfe00;
			16'hd057: y = 16'hfe00;
			16'hd058: y = 16'hfe00;
			16'hd059: y = 16'hfe00;
			16'hd05a: y = 16'hfe00;
			16'hd05b: y = 16'hfe00;
			16'hd05c: y = 16'hfe00;
			16'hd05d: y = 16'hfe00;
			16'hd05e: y = 16'hfe00;
			16'hd05f: y = 16'hfe00;
			16'hd060: y = 16'hfe00;
			16'hd061: y = 16'hfe00;
			16'hd062: y = 16'hfe00;
			16'hd063: y = 16'hfe00;
			16'hd064: y = 16'hfe00;
			16'hd065: y = 16'hfe00;
			16'hd066: y = 16'hfe00;
			16'hd067: y = 16'hfe00;
			16'hd068: y = 16'hfe00;
			16'hd069: y = 16'hfe00;
			16'hd06a: y = 16'hfe00;
			16'hd06b: y = 16'hfe00;
			16'hd06c: y = 16'hfe00;
			16'hd06d: y = 16'hfe00;
			16'hd06e: y = 16'hfe00;
			16'hd06f: y = 16'hfe00;
			16'hd070: y = 16'hfe00;
			16'hd071: y = 16'hfe00;
			16'hd072: y = 16'hfe00;
			16'hd073: y = 16'hfe00;
			16'hd074: y = 16'hfe00;
			16'hd075: y = 16'hfe00;
			16'hd076: y = 16'hfe00;
			16'hd077: y = 16'hfe00;
			16'hd078: y = 16'hfe00;
			16'hd079: y = 16'hfe00;
			16'hd07a: y = 16'hfe00;
			16'hd07b: y = 16'hfe00;
			16'hd07c: y = 16'hfe00;
			16'hd07d: y = 16'hfe00;
			16'hd07e: y = 16'hfe00;
			16'hd07f: y = 16'hfe00;
			16'hd080: y = 16'hfe00;
			16'hd081: y = 16'hfe00;
			16'hd082: y = 16'hfe00;
			16'hd083: y = 16'hfe00;
			16'hd084: y = 16'hfe00;
			16'hd085: y = 16'hfe00;
			16'hd086: y = 16'hfe00;
			16'hd087: y = 16'hfe00;
			16'hd088: y = 16'hfe00;
			16'hd089: y = 16'hfe00;
			16'hd08a: y = 16'hfe00;
			16'hd08b: y = 16'hfe00;
			16'hd08c: y = 16'hfe00;
			16'hd08d: y = 16'hfe00;
			16'hd08e: y = 16'hfe00;
			16'hd08f: y = 16'hfe00;
			16'hd090: y = 16'hfe00;
			16'hd091: y = 16'hfe00;
			16'hd092: y = 16'hfe00;
			16'hd093: y = 16'hfe00;
			16'hd094: y = 16'hfe00;
			16'hd095: y = 16'hfe00;
			16'hd096: y = 16'hfe00;
			16'hd097: y = 16'hfe00;
			16'hd098: y = 16'hfe00;
			16'hd099: y = 16'hfe00;
			16'hd09a: y = 16'hfe00;
			16'hd09b: y = 16'hfe00;
			16'hd09c: y = 16'hfe00;
			16'hd09d: y = 16'hfe00;
			16'hd09e: y = 16'hfe00;
			16'hd09f: y = 16'hfe00;
			16'hd0a0: y = 16'hfe00;
			16'hd0a1: y = 16'hfe00;
			16'hd0a2: y = 16'hfe00;
			16'hd0a3: y = 16'hfe00;
			16'hd0a4: y = 16'hfe00;
			16'hd0a5: y = 16'hfe00;
			16'hd0a6: y = 16'hfe00;
			16'hd0a7: y = 16'hfe00;
			16'hd0a8: y = 16'hfe00;
			16'hd0a9: y = 16'hfe00;
			16'hd0aa: y = 16'hfe00;
			16'hd0ab: y = 16'hfe00;
			16'hd0ac: y = 16'hfe00;
			16'hd0ad: y = 16'hfe00;
			16'hd0ae: y = 16'hfe00;
			16'hd0af: y = 16'hfe00;
			16'hd0b0: y = 16'hfe00;
			16'hd0b1: y = 16'hfe00;
			16'hd0b2: y = 16'hfe00;
			16'hd0b3: y = 16'hfe00;
			16'hd0b4: y = 16'hfe00;
			16'hd0b5: y = 16'hfe00;
			16'hd0b6: y = 16'hfe00;
			16'hd0b7: y = 16'hfe00;
			16'hd0b8: y = 16'hfe00;
			16'hd0b9: y = 16'hfe00;
			16'hd0ba: y = 16'hfe00;
			16'hd0bb: y = 16'hfe00;
			16'hd0bc: y = 16'hfe00;
			16'hd0bd: y = 16'hfe00;
			16'hd0be: y = 16'hfe00;
			16'hd0bf: y = 16'hfe00;
			16'hd0c0: y = 16'hfe00;
			16'hd0c1: y = 16'hfe00;
			16'hd0c2: y = 16'hfe00;
			16'hd0c3: y = 16'hfe00;
			16'hd0c4: y = 16'hfe00;
			16'hd0c5: y = 16'hfe00;
			16'hd0c6: y = 16'hfe00;
			16'hd0c7: y = 16'hfe00;
			16'hd0c8: y = 16'hfe00;
			16'hd0c9: y = 16'hfe00;
			16'hd0ca: y = 16'hfe00;
			16'hd0cb: y = 16'hfe00;
			16'hd0cc: y = 16'hfe00;
			16'hd0cd: y = 16'hfe00;
			16'hd0ce: y = 16'hfe00;
			16'hd0cf: y = 16'hfe00;
			16'hd0d0: y = 16'hfe00;
			16'hd0d1: y = 16'hfe00;
			16'hd0d2: y = 16'hfe00;
			16'hd0d3: y = 16'hfe00;
			16'hd0d4: y = 16'hfe00;
			16'hd0d5: y = 16'hfe00;
			16'hd0d6: y = 16'hfe00;
			16'hd0d7: y = 16'hfe00;
			16'hd0d8: y = 16'hfe00;
			16'hd0d9: y = 16'hfe00;
			16'hd0da: y = 16'hfe00;
			16'hd0db: y = 16'hfe00;
			16'hd0dc: y = 16'hfe00;
			16'hd0dd: y = 16'hfe00;
			16'hd0de: y = 16'hfe00;
			16'hd0df: y = 16'hfe00;
			16'hd0e0: y = 16'hfe00;
			16'hd0e1: y = 16'hfe00;
			16'hd0e2: y = 16'hfe00;
			16'hd0e3: y = 16'hfe00;
			16'hd0e4: y = 16'hfe00;
			16'hd0e5: y = 16'hfe00;
			16'hd0e6: y = 16'hfe00;
			16'hd0e7: y = 16'hfe00;
			16'hd0e8: y = 16'hfe00;
			16'hd0e9: y = 16'hfe00;
			16'hd0ea: y = 16'hfe00;
			16'hd0eb: y = 16'hfe00;
			16'hd0ec: y = 16'hfe00;
			16'hd0ed: y = 16'hfe00;
			16'hd0ee: y = 16'hfe00;
			16'hd0ef: y = 16'hfe00;
			16'hd0f0: y = 16'hfe00;
			16'hd0f1: y = 16'hfe00;
			16'hd0f2: y = 16'hfe00;
			16'hd0f3: y = 16'hfe00;
			16'hd0f4: y = 16'hfe00;
			16'hd0f5: y = 16'hfe00;
			16'hd0f6: y = 16'hfe00;
			16'hd0f7: y = 16'hfe00;
			16'hd0f8: y = 16'hfe00;
			16'hd0f9: y = 16'hfe00;
			16'hd0fa: y = 16'hfe00;
			16'hd0fb: y = 16'hfe00;
			16'hd0fc: y = 16'hfe00;
			16'hd0fd: y = 16'hfe00;
			16'hd0fe: y = 16'hfe00;
			16'hd0ff: y = 16'hfe00;
			16'hd100: y = 16'hfe00;
			16'hd101: y = 16'hfe00;
			16'hd102: y = 16'hfe00;
			16'hd103: y = 16'hfe00;
			16'hd104: y = 16'hfe00;
			16'hd105: y = 16'hfe00;
			16'hd106: y = 16'hfe00;
			16'hd107: y = 16'hfe00;
			16'hd108: y = 16'hfe00;
			16'hd109: y = 16'hfe00;
			16'hd10a: y = 16'hfe00;
			16'hd10b: y = 16'hfe00;
			16'hd10c: y = 16'hfe00;
			16'hd10d: y = 16'hfe00;
			16'hd10e: y = 16'hfe00;
			16'hd10f: y = 16'hfe00;
			16'hd110: y = 16'hfe00;
			16'hd111: y = 16'hfe00;
			16'hd112: y = 16'hfe00;
			16'hd113: y = 16'hfe00;
			16'hd114: y = 16'hfe00;
			16'hd115: y = 16'hfe00;
			16'hd116: y = 16'hfe00;
			16'hd117: y = 16'hfe00;
			16'hd118: y = 16'hfe00;
			16'hd119: y = 16'hfe00;
			16'hd11a: y = 16'hfe00;
			16'hd11b: y = 16'hfe00;
			16'hd11c: y = 16'hfe00;
			16'hd11d: y = 16'hfe00;
			16'hd11e: y = 16'hfe00;
			16'hd11f: y = 16'hfe00;
			16'hd120: y = 16'hfe00;
			16'hd121: y = 16'hfe00;
			16'hd122: y = 16'hfe00;
			16'hd123: y = 16'hfe00;
			16'hd124: y = 16'hfe00;
			16'hd125: y = 16'hfe00;
			16'hd126: y = 16'hfe00;
			16'hd127: y = 16'hfe00;
			16'hd128: y = 16'hfe00;
			16'hd129: y = 16'hfe00;
			16'hd12a: y = 16'hfe00;
			16'hd12b: y = 16'hfe00;
			16'hd12c: y = 16'hfe00;
			16'hd12d: y = 16'hfe00;
			16'hd12e: y = 16'hfe00;
			16'hd12f: y = 16'hfe00;
			16'hd130: y = 16'hfe00;
			16'hd131: y = 16'hfe00;
			16'hd132: y = 16'hfe00;
			16'hd133: y = 16'hfe00;
			16'hd134: y = 16'hfe00;
			16'hd135: y = 16'hfe00;
			16'hd136: y = 16'hfe00;
			16'hd137: y = 16'hfe00;
			16'hd138: y = 16'hfe00;
			16'hd139: y = 16'hfe00;
			16'hd13a: y = 16'hfe00;
			16'hd13b: y = 16'hfe00;
			16'hd13c: y = 16'hfe00;
			16'hd13d: y = 16'hfe00;
			16'hd13e: y = 16'hfe00;
			16'hd13f: y = 16'hfe00;
			16'hd140: y = 16'hfe00;
			16'hd141: y = 16'hfe00;
			16'hd142: y = 16'hfe00;
			16'hd143: y = 16'hfe00;
			16'hd144: y = 16'hfe00;
			16'hd145: y = 16'hfe00;
			16'hd146: y = 16'hfe00;
			16'hd147: y = 16'hfe00;
			16'hd148: y = 16'hfe00;
			16'hd149: y = 16'hfe00;
			16'hd14a: y = 16'hfe00;
			16'hd14b: y = 16'hfe00;
			16'hd14c: y = 16'hfe00;
			16'hd14d: y = 16'hfe00;
			16'hd14e: y = 16'hfe00;
			16'hd14f: y = 16'hfe00;
			16'hd150: y = 16'hfe00;
			16'hd151: y = 16'hfe00;
			16'hd152: y = 16'hfe00;
			16'hd153: y = 16'hfe00;
			16'hd154: y = 16'hfe00;
			16'hd155: y = 16'hfe00;
			16'hd156: y = 16'hfe00;
			16'hd157: y = 16'hfe00;
			16'hd158: y = 16'hfe00;
			16'hd159: y = 16'hfe00;
			16'hd15a: y = 16'hfe00;
			16'hd15b: y = 16'hfe00;
			16'hd15c: y = 16'hfe00;
			16'hd15d: y = 16'hfe00;
			16'hd15e: y = 16'hfe00;
			16'hd15f: y = 16'hfe00;
			16'hd160: y = 16'hfe00;
			16'hd161: y = 16'hfe00;
			16'hd162: y = 16'hfe00;
			16'hd163: y = 16'hfe00;
			16'hd164: y = 16'hfe00;
			16'hd165: y = 16'hfe00;
			16'hd166: y = 16'hfe00;
			16'hd167: y = 16'hfe00;
			16'hd168: y = 16'hfe00;
			16'hd169: y = 16'hfe00;
			16'hd16a: y = 16'hfe00;
			16'hd16b: y = 16'hfe00;
			16'hd16c: y = 16'hfe00;
			16'hd16d: y = 16'hfe00;
			16'hd16e: y = 16'hfe00;
			16'hd16f: y = 16'hfe00;
			16'hd170: y = 16'hfe00;
			16'hd171: y = 16'hfe00;
			16'hd172: y = 16'hfe00;
			16'hd173: y = 16'hfe00;
			16'hd174: y = 16'hfe00;
			16'hd175: y = 16'hfe00;
			16'hd176: y = 16'hfe00;
			16'hd177: y = 16'hfe00;
			16'hd178: y = 16'hfe00;
			16'hd179: y = 16'hfe00;
			16'hd17a: y = 16'hfe00;
			16'hd17b: y = 16'hfe00;
			16'hd17c: y = 16'hfe00;
			16'hd17d: y = 16'hfe00;
			16'hd17e: y = 16'hfe00;
			16'hd17f: y = 16'hfe00;
			16'hd180: y = 16'hfe00;
			16'hd181: y = 16'hfe00;
			16'hd182: y = 16'hfe00;
			16'hd183: y = 16'hfe00;
			16'hd184: y = 16'hfe00;
			16'hd185: y = 16'hfe00;
			16'hd186: y = 16'hfe00;
			16'hd187: y = 16'hfe00;
			16'hd188: y = 16'hfe00;
			16'hd189: y = 16'hfe00;
			16'hd18a: y = 16'hfe00;
			16'hd18b: y = 16'hfe00;
			16'hd18c: y = 16'hfe00;
			16'hd18d: y = 16'hfe00;
			16'hd18e: y = 16'hfe00;
			16'hd18f: y = 16'hfe00;
			16'hd190: y = 16'hfe00;
			16'hd191: y = 16'hfe00;
			16'hd192: y = 16'hfe00;
			16'hd193: y = 16'hfe00;
			16'hd194: y = 16'hfe00;
			16'hd195: y = 16'hfe00;
			16'hd196: y = 16'hfe00;
			16'hd197: y = 16'hfe00;
			16'hd198: y = 16'hfe00;
			16'hd199: y = 16'hfe00;
			16'hd19a: y = 16'hfe00;
			16'hd19b: y = 16'hfe00;
			16'hd19c: y = 16'hfe00;
			16'hd19d: y = 16'hfe00;
			16'hd19e: y = 16'hfe00;
			16'hd19f: y = 16'hfe00;
			16'hd1a0: y = 16'hfe00;
			16'hd1a1: y = 16'hfe00;
			16'hd1a2: y = 16'hfe00;
			16'hd1a3: y = 16'hfe00;
			16'hd1a4: y = 16'hfe00;
			16'hd1a5: y = 16'hfe00;
			16'hd1a6: y = 16'hfe00;
			16'hd1a7: y = 16'hfe00;
			16'hd1a8: y = 16'hfe00;
			16'hd1a9: y = 16'hfe00;
			16'hd1aa: y = 16'hfe00;
			16'hd1ab: y = 16'hfe00;
			16'hd1ac: y = 16'hfe00;
			16'hd1ad: y = 16'hfe00;
			16'hd1ae: y = 16'hfe00;
			16'hd1af: y = 16'hfe00;
			16'hd1b0: y = 16'hfe00;
			16'hd1b1: y = 16'hfe00;
			16'hd1b2: y = 16'hfe00;
			16'hd1b3: y = 16'hfe00;
			16'hd1b4: y = 16'hfe00;
			16'hd1b5: y = 16'hfe00;
			16'hd1b6: y = 16'hfe00;
			16'hd1b7: y = 16'hfe00;
			16'hd1b8: y = 16'hfe00;
			16'hd1b9: y = 16'hfe00;
			16'hd1ba: y = 16'hfe00;
			16'hd1bb: y = 16'hfe00;
			16'hd1bc: y = 16'hfe00;
			16'hd1bd: y = 16'hfe00;
			16'hd1be: y = 16'hfe00;
			16'hd1bf: y = 16'hfe00;
			16'hd1c0: y = 16'hfe00;
			16'hd1c1: y = 16'hfe00;
			16'hd1c2: y = 16'hfe00;
			16'hd1c3: y = 16'hfe00;
			16'hd1c4: y = 16'hfe00;
			16'hd1c5: y = 16'hfe00;
			16'hd1c6: y = 16'hfe00;
			16'hd1c7: y = 16'hfe00;
			16'hd1c8: y = 16'hfe00;
			16'hd1c9: y = 16'hfe00;
			16'hd1ca: y = 16'hfe00;
			16'hd1cb: y = 16'hfe00;
			16'hd1cc: y = 16'hfe00;
			16'hd1cd: y = 16'hfe00;
			16'hd1ce: y = 16'hfe00;
			16'hd1cf: y = 16'hfe00;
			16'hd1d0: y = 16'hfe00;
			16'hd1d1: y = 16'hfe00;
			16'hd1d2: y = 16'hfe00;
			16'hd1d3: y = 16'hfe00;
			16'hd1d4: y = 16'hfe00;
			16'hd1d5: y = 16'hfe00;
			16'hd1d6: y = 16'hfe00;
			16'hd1d7: y = 16'hfe00;
			16'hd1d8: y = 16'hfe00;
			16'hd1d9: y = 16'hfe00;
			16'hd1da: y = 16'hfe00;
			16'hd1db: y = 16'hfe00;
			16'hd1dc: y = 16'hfe00;
			16'hd1dd: y = 16'hfe00;
			16'hd1de: y = 16'hfe00;
			16'hd1df: y = 16'hfe00;
			16'hd1e0: y = 16'hfe00;
			16'hd1e1: y = 16'hfe00;
			16'hd1e2: y = 16'hfe00;
			16'hd1e3: y = 16'hfe00;
			16'hd1e4: y = 16'hfe00;
			16'hd1e5: y = 16'hfe00;
			16'hd1e6: y = 16'hfe00;
			16'hd1e7: y = 16'hfe00;
			16'hd1e8: y = 16'hfe00;
			16'hd1e9: y = 16'hfe00;
			16'hd1ea: y = 16'hfe00;
			16'hd1eb: y = 16'hfe00;
			16'hd1ec: y = 16'hfe00;
			16'hd1ed: y = 16'hfe00;
			16'hd1ee: y = 16'hfe00;
			16'hd1ef: y = 16'hfe00;
			16'hd1f0: y = 16'hfe00;
			16'hd1f1: y = 16'hfe00;
			16'hd1f2: y = 16'hfe00;
			16'hd1f3: y = 16'hfe00;
			16'hd1f4: y = 16'hfe00;
			16'hd1f5: y = 16'hfe00;
			16'hd1f6: y = 16'hfe00;
			16'hd1f7: y = 16'hfe00;
			16'hd1f8: y = 16'hfe00;
			16'hd1f9: y = 16'hfe00;
			16'hd1fa: y = 16'hfe00;
			16'hd1fb: y = 16'hfe00;
			16'hd1fc: y = 16'hfe00;
			16'hd1fd: y = 16'hfe00;
			16'hd1fe: y = 16'hfe00;
			16'hd1ff: y = 16'hfe00;
			16'hd200: y = 16'hfe00;
			16'hd201: y = 16'hfe00;
			16'hd202: y = 16'hfe00;
			16'hd203: y = 16'hfe00;
			16'hd204: y = 16'hfe00;
			16'hd205: y = 16'hfe00;
			16'hd206: y = 16'hfe00;
			16'hd207: y = 16'hfe00;
			16'hd208: y = 16'hfe00;
			16'hd209: y = 16'hfe00;
			16'hd20a: y = 16'hfe00;
			16'hd20b: y = 16'hfe00;
			16'hd20c: y = 16'hfe00;
			16'hd20d: y = 16'hfe00;
			16'hd20e: y = 16'hfe00;
			16'hd20f: y = 16'hfe00;
			16'hd210: y = 16'hfe00;
			16'hd211: y = 16'hfe00;
			16'hd212: y = 16'hfe00;
			16'hd213: y = 16'hfe00;
			16'hd214: y = 16'hfe00;
			16'hd215: y = 16'hfe00;
			16'hd216: y = 16'hfe00;
			16'hd217: y = 16'hfe00;
			16'hd218: y = 16'hfe00;
			16'hd219: y = 16'hfe00;
			16'hd21a: y = 16'hfe00;
			16'hd21b: y = 16'hfe00;
			16'hd21c: y = 16'hfe00;
			16'hd21d: y = 16'hfe00;
			16'hd21e: y = 16'hfe00;
			16'hd21f: y = 16'hfe00;
			16'hd220: y = 16'hfe00;
			16'hd221: y = 16'hfe00;
			16'hd222: y = 16'hfe00;
			16'hd223: y = 16'hfe00;
			16'hd224: y = 16'hfe00;
			16'hd225: y = 16'hfe00;
			16'hd226: y = 16'hfe00;
			16'hd227: y = 16'hfe00;
			16'hd228: y = 16'hfe00;
			16'hd229: y = 16'hfe00;
			16'hd22a: y = 16'hfe00;
			16'hd22b: y = 16'hfe00;
			16'hd22c: y = 16'hfe00;
			16'hd22d: y = 16'hfe00;
			16'hd22e: y = 16'hfe00;
			16'hd22f: y = 16'hfe00;
			16'hd230: y = 16'hfe00;
			16'hd231: y = 16'hfe00;
			16'hd232: y = 16'hfe00;
			16'hd233: y = 16'hfe00;
			16'hd234: y = 16'hfe00;
			16'hd235: y = 16'hfe00;
			16'hd236: y = 16'hfe00;
			16'hd237: y = 16'hfe00;
			16'hd238: y = 16'hfe00;
			16'hd239: y = 16'hfe00;
			16'hd23a: y = 16'hfe00;
			16'hd23b: y = 16'hfe00;
			16'hd23c: y = 16'hfe00;
			16'hd23d: y = 16'hfe00;
			16'hd23e: y = 16'hfe00;
			16'hd23f: y = 16'hfe00;
			16'hd240: y = 16'hfe00;
			16'hd241: y = 16'hfe00;
			16'hd242: y = 16'hfe00;
			16'hd243: y = 16'hfe00;
			16'hd244: y = 16'hfe00;
			16'hd245: y = 16'hfe00;
			16'hd246: y = 16'hfe00;
			16'hd247: y = 16'hfe00;
			16'hd248: y = 16'hfe00;
			16'hd249: y = 16'hfe00;
			16'hd24a: y = 16'hfe00;
			16'hd24b: y = 16'hfe00;
			16'hd24c: y = 16'hfe00;
			16'hd24d: y = 16'hfe00;
			16'hd24e: y = 16'hfe00;
			16'hd24f: y = 16'hfe00;
			16'hd250: y = 16'hfe00;
			16'hd251: y = 16'hfe00;
			16'hd252: y = 16'hfe00;
			16'hd253: y = 16'hfe00;
			16'hd254: y = 16'hfe00;
			16'hd255: y = 16'hfe00;
			16'hd256: y = 16'hfe00;
			16'hd257: y = 16'hfe00;
			16'hd258: y = 16'hfe00;
			16'hd259: y = 16'hfe00;
			16'hd25a: y = 16'hfe00;
			16'hd25b: y = 16'hfe00;
			16'hd25c: y = 16'hfe00;
			16'hd25d: y = 16'hfe00;
			16'hd25e: y = 16'hfe00;
			16'hd25f: y = 16'hfe00;
			16'hd260: y = 16'hfe00;
			16'hd261: y = 16'hfe00;
			16'hd262: y = 16'hfe00;
			16'hd263: y = 16'hfe00;
			16'hd264: y = 16'hfe00;
			16'hd265: y = 16'hfe00;
			16'hd266: y = 16'hfe00;
			16'hd267: y = 16'hfe00;
			16'hd268: y = 16'hfe00;
			16'hd269: y = 16'hfe00;
			16'hd26a: y = 16'hfe00;
			16'hd26b: y = 16'hfe00;
			16'hd26c: y = 16'hfe00;
			16'hd26d: y = 16'hfe00;
			16'hd26e: y = 16'hfe00;
			16'hd26f: y = 16'hfe00;
			16'hd270: y = 16'hfe00;
			16'hd271: y = 16'hfe00;
			16'hd272: y = 16'hfe00;
			16'hd273: y = 16'hfe00;
			16'hd274: y = 16'hfe00;
			16'hd275: y = 16'hfe00;
			16'hd276: y = 16'hfe00;
			16'hd277: y = 16'hfe00;
			16'hd278: y = 16'hfe00;
			16'hd279: y = 16'hfe00;
			16'hd27a: y = 16'hfe00;
			16'hd27b: y = 16'hfe00;
			16'hd27c: y = 16'hfe00;
			16'hd27d: y = 16'hfe00;
			16'hd27e: y = 16'hfe00;
			16'hd27f: y = 16'hfe00;
			16'hd280: y = 16'hfe00;
			16'hd281: y = 16'hfe00;
			16'hd282: y = 16'hfe00;
			16'hd283: y = 16'hfe00;
			16'hd284: y = 16'hfe00;
			16'hd285: y = 16'hfe00;
			16'hd286: y = 16'hfe00;
			16'hd287: y = 16'hfe00;
			16'hd288: y = 16'hfe00;
			16'hd289: y = 16'hfe00;
			16'hd28a: y = 16'hfe00;
			16'hd28b: y = 16'hfe00;
			16'hd28c: y = 16'hfe00;
			16'hd28d: y = 16'hfe00;
			16'hd28e: y = 16'hfe00;
			16'hd28f: y = 16'hfe00;
			16'hd290: y = 16'hfe00;
			16'hd291: y = 16'hfe00;
			16'hd292: y = 16'hfe00;
			16'hd293: y = 16'hfe00;
			16'hd294: y = 16'hfe00;
			16'hd295: y = 16'hfe00;
			16'hd296: y = 16'hfe00;
			16'hd297: y = 16'hfe00;
			16'hd298: y = 16'hfe00;
			16'hd299: y = 16'hfe00;
			16'hd29a: y = 16'hfe00;
			16'hd29b: y = 16'hfe00;
			16'hd29c: y = 16'hfe00;
			16'hd29d: y = 16'hfe00;
			16'hd29e: y = 16'hfe00;
			16'hd29f: y = 16'hfe00;
			16'hd2a0: y = 16'hfe00;
			16'hd2a1: y = 16'hfe00;
			16'hd2a2: y = 16'hfe00;
			16'hd2a3: y = 16'hfe00;
			16'hd2a4: y = 16'hfe00;
			16'hd2a5: y = 16'hfe00;
			16'hd2a6: y = 16'hfe00;
			16'hd2a7: y = 16'hfe00;
			16'hd2a8: y = 16'hfe00;
			16'hd2a9: y = 16'hfe00;
			16'hd2aa: y = 16'hfe00;
			16'hd2ab: y = 16'hfe00;
			16'hd2ac: y = 16'hfe00;
			16'hd2ad: y = 16'hfe00;
			16'hd2ae: y = 16'hfe00;
			16'hd2af: y = 16'hfe00;
			16'hd2b0: y = 16'hfe00;
			16'hd2b1: y = 16'hfe00;
			16'hd2b2: y = 16'hfe00;
			16'hd2b3: y = 16'hfe00;
			16'hd2b4: y = 16'hfe00;
			16'hd2b5: y = 16'hfe00;
			16'hd2b6: y = 16'hfe00;
			16'hd2b7: y = 16'hfe00;
			16'hd2b8: y = 16'hfe00;
			16'hd2b9: y = 16'hfe00;
			16'hd2ba: y = 16'hfe00;
			16'hd2bb: y = 16'hfe00;
			16'hd2bc: y = 16'hfe00;
			16'hd2bd: y = 16'hfe00;
			16'hd2be: y = 16'hfe00;
			16'hd2bf: y = 16'hfe00;
			16'hd2c0: y = 16'hfe00;
			16'hd2c1: y = 16'hfe00;
			16'hd2c2: y = 16'hfe00;
			16'hd2c3: y = 16'hfe00;
			16'hd2c4: y = 16'hfe00;
			16'hd2c5: y = 16'hfe00;
			16'hd2c6: y = 16'hfe00;
			16'hd2c7: y = 16'hfe00;
			16'hd2c8: y = 16'hfe00;
			16'hd2c9: y = 16'hfe00;
			16'hd2ca: y = 16'hfe00;
			16'hd2cb: y = 16'hfe00;
			16'hd2cc: y = 16'hfe00;
			16'hd2cd: y = 16'hfe00;
			16'hd2ce: y = 16'hfe00;
			16'hd2cf: y = 16'hfe00;
			16'hd2d0: y = 16'hfe00;
			16'hd2d1: y = 16'hfe00;
			16'hd2d2: y = 16'hfe00;
			16'hd2d3: y = 16'hfe00;
			16'hd2d4: y = 16'hfe00;
			16'hd2d5: y = 16'hfe00;
			16'hd2d6: y = 16'hfe00;
			16'hd2d7: y = 16'hfe00;
			16'hd2d8: y = 16'hfe00;
			16'hd2d9: y = 16'hfe00;
			16'hd2da: y = 16'hfe00;
			16'hd2db: y = 16'hfe00;
			16'hd2dc: y = 16'hfe00;
			16'hd2dd: y = 16'hfe00;
			16'hd2de: y = 16'hfe00;
			16'hd2df: y = 16'hfe00;
			16'hd2e0: y = 16'hfe00;
			16'hd2e1: y = 16'hfe00;
			16'hd2e2: y = 16'hfe00;
			16'hd2e3: y = 16'hfe00;
			16'hd2e4: y = 16'hfe00;
			16'hd2e5: y = 16'hfe00;
			16'hd2e6: y = 16'hfe00;
			16'hd2e7: y = 16'hfe00;
			16'hd2e8: y = 16'hfe00;
			16'hd2e9: y = 16'hfe00;
			16'hd2ea: y = 16'hfe00;
			16'hd2eb: y = 16'hfe00;
			16'hd2ec: y = 16'hfe00;
			16'hd2ed: y = 16'hfe00;
			16'hd2ee: y = 16'hfe00;
			16'hd2ef: y = 16'hfe00;
			16'hd2f0: y = 16'hfe00;
			16'hd2f1: y = 16'hfe00;
			16'hd2f2: y = 16'hfe00;
			16'hd2f3: y = 16'hfe00;
			16'hd2f4: y = 16'hfe00;
			16'hd2f5: y = 16'hfe00;
			16'hd2f6: y = 16'hfe00;
			16'hd2f7: y = 16'hfe00;
			16'hd2f8: y = 16'hfe00;
			16'hd2f9: y = 16'hfe00;
			16'hd2fa: y = 16'hfe00;
			16'hd2fb: y = 16'hfe00;
			16'hd2fc: y = 16'hfe00;
			16'hd2fd: y = 16'hfe00;
			16'hd2fe: y = 16'hfe00;
			16'hd2ff: y = 16'hfe00;
			16'hd300: y = 16'hfe00;
			16'hd301: y = 16'hfe00;
			16'hd302: y = 16'hfe00;
			16'hd303: y = 16'hfe00;
			16'hd304: y = 16'hfe00;
			16'hd305: y = 16'hfe00;
			16'hd306: y = 16'hfe00;
			16'hd307: y = 16'hfe00;
			16'hd308: y = 16'hfe00;
			16'hd309: y = 16'hfe00;
			16'hd30a: y = 16'hfe00;
			16'hd30b: y = 16'hfe00;
			16'hd30c: y = 16'hfe00;
			16'hd30d: y = 16'hfe00;
			16'hd30e: y = 16'hfe00;
			16'hd30f: y = 16'hfe00;
			16'hd310: y = 16'hfe00;
			16'hd311: y = 16'hfe00;
			16'hd312: y = 16'hfe00;
			16'hd313: y = 16'hfe00;
			16'hd314: y = 16'hfe00;
			16'hd315: y = 16'hfe00;
			16'hd316: y = 16'hfe00;
			16'hd317: y = 16'hfe00;
			16'hd318: y = 16'hfe00;
			16'hd319: y = 16'hfe00;
			16'hd31a: y = 16'hfe00;
			16'hd31b: y = 16'hfe00;
			16'hd31c: y = 16'hfe00;
			16'hd31d: y = 16'hfe00;
			16'hd31e: y = 16'hfe00;
			16'hd31f: y = 16'hfe00;
			16'hd320: y = 16'hfe00;
			16'hd321: y = 16'hfe00;
			16'hd322: y = 16'hfe00;
			16'hd323: y = 16'hfe00;
			16'hd324: y = 16'hfe00;
			16'hd325: y = 16'hfe00;
			16'hd326: y = 16'hfe00;
			16'hd327: y = 16'hfe00;
			16'hd328: y = 16'hfe00;
			16'hd329: y = 16'hfe00;
			16'hd32a: y = 16'hfe00;
			16'hd32b: y = 16'hfe00;
			16'hd32c: y = 16'hfe00;
			16'hd32d: y = 16'hfe00;
			16'hd32e: y = 16'hfe00;
			16'hd32f: y = 16'hfe00;
			16'hd330: y = 16'hfe00;
			16'hd331: y = 16'hfe00;
			16'hd332: y = 16'hfe00;
			16'hd333: y = 16'hfe00;
			16'hd334: y = 16'hfe00;
			16'hd335: y = 16'hfe00;
			16'hd336: y = 16'hfe00;
			16'hd337: y = 16'hfe00;
			16'hd338: y = 16'hfe00;
			16'hd339: y = 16'hfe00;
			16'hd33a: y = 16'hfe00;
			16'hd33b: y = 16'hfe00;
			16'hd33c: y = 16'hfe00;
			16'hd33d: y = 16'hfe00;
			16'hd33e: y = 16'hfe00;
			16'hd33f: y = 16'hfe00;
			16'hd340: y = 16'hfe00;
			16'hd341: y = 16'hfe00;
			16'hd342: y = 16'hfe00;
			16'hd343: y = 16'hfe00;
			16'hd344: y = 16'hfe00;
			16'hd345: y = 16'hfe00;
			16'hd346: y = 16'hfe00;
			16'hd347: y = 16'hfe00;
			16'hd348: y = 16'hfe00;
			16'hd349: y = 16'hfe00;
			16'hd34a: y = 16'hfe00;
			16'hd34b: y = 16'hfe00;
			16'hd34c: y = 16'hfe00;
			16'hd34d: y = 16'hfe00;
			16'hd34e: y = 16'hfe00;
			16'hd34f: y = 16'hfe00;
			16'hd350: y = 16'hfe00;
			16'hd351: y = 16'hfe00;
			16'hd352: y = 16'hfe00;
			16'hd353: y = 16'hfe00;
			16'hd354: y = 16'hfe00;
			16'hd355: y = 16'hfe00;
			16'hd356: y = 16'hfe00;
			16'hd357: y = 16'hfe00;
			16'hd358: y = 16'hfe00;
			16'hd359: y = 16'hfe00;
			16'hd35a: y = 16'hfe00;
			16'hd35b: y = 16'hfe00;
			16'hd35c: y = 16'hfe00;
			16'hd35d: y = 16'hfe00;
			16'hd35e: y = 16'hfe00;
			16'hd35f: y = 16'hfe00;
			16'hd360: y = 16'hfe00;
			16'hd361: y = 16'hfe00;
			16'hd362: y = 16'hfe00;
			16'hd363: y = 16'hfe00;
			16'hd364: y = 16'hfe00;
			16'hd365: y = 16'hfe00;
			16'hd366: y = 16'hfe00;
			16'hd367: y = 16'hfe00;
			16'hd368: y = 16'hfe00;
			16'hd369: y = 16'hfe00;
			16'hd36a: y = 16'hfe00;
			16'hd36b: y = 16'hfe00;
			16'hd36c: y = 16'hfe00;
			16'hd36d: y = 16'hfe00;
			16'hd36e: y = 16'hfe00;
			16'hd36f: y = 16'hfe00;
			16'hd370: y = 16'hfe00;
			16'hd371: y = 16'hfe00;
			16'hd372: y = 16'hfe00;
			16'hd373: y = 16'hfe00;
			16'hd374: y = 16'hfe00;
			16'hd375: y = 16'hfe00;
			16'hd376: y = 16'hfe00;
			16'hd377: y = 16'hfe00;
			16'hd378: y = 16'hfe00;
			16'hd379: y = 16'hfe00;
			16'hd37a: y = 16'hfe00;
			16'hd37b: y = 16'hfe00;
			16'hd37c: y = 16'hfe00;
			16'hd37d: y = 16'hfe00;
			16'hd37e: y = 16'hfe00;
			16'hd37f: y = 16'hfe00;
			16'hd380: y = 16'hfe00;
			16'hd381: y = 16'hfe00;
			16'hd382: y = 16'hfe00;
			16'hd383: y = 16'hfe00;
			16'hd384: y = 16'hfe00;
			16'hd385: y = 16'hfe00;
			16'hd386: y = 16'hfe00;
			16'hd387: y = 16'hfe00;
			16'hd388: y = 16'hfe00;
			16'hd389: y = 16'hfe00;
			16'hd38a: y = 16'hfe00;
			16'hd38b: y = 16'hfe00;
			16'hd38c: y = 16'hfe00;
			16'hd38d: y = 16'hfe00;
			16'hd38e: y = 16'hfe00;
			16'hd38f: y = 16'hfe00;
			16'hd390: y = 16'hfe00;
			16'hd391: y = 16'hfe00;
			16'hd392: y = 16'hfe00;
			16'hd393: y = 16'hfe00;
			16'hd394: y = 16'hfe00;
			16'hd395: y = 16'hfe00;
			16'hd396: y = 16'hfe00;
			16'hd397: y = 16'hfe00;
			16'hd398: y = 16'hfe00;
			16'hd399: y = 16'hfe00;
			16'hd39a: y = 16'hfe00;
			16'hd39b: y = 16'hfe00;
			16'hd39c: y = 16'hfe00;
			16'hd39d: y = 16'hfe00;
			16'hd39e: y = 16'hfe00;
			16'hd39f: y = 16'hfe00;
			16'hd3a0: y = 16'hfe00;
			16'hd3a1: y = 16'hfe00;
			16'hd3a2: y = 16'hfe00;
			16'hd3a3: y = 16'hfe00;
			16'hd3a4: y = 16'hfe00;
			16'hd3a5: y = 16'hfe00;
			16'hd3a6: y = 16'hfe00;
			16'hd3a7: y = 16'hfe00;
			16'hd3a8: y = 16'hfe00;
			16'hd3a9: y = 16'hfe00;
			16'hd3aa: y = 16'hfe00;
			16'hd3ab: y = 16'hfe00;
			16'hd3ac: y = 16'hfe00;
			16'hd3ad: y = 16'hfe00;
			16'hd3ae: y = 16'hfe00;
			16'hd3af: y = 16'hfe00;
			16'hd3b0: y = 16'hfe00;
			16'hd3b1: y = 16'hfe00;
			16'hd3b2: y = 16'hfe00;
			16'hd3b3: y = 16'hfe00;
			16'hd3b4: y = 16'hfe00;
			16'hd3b5: y = 16'hfe00;
			16'hd3b6: y = 16'hfe00;
			16'hd3b7: y = 16'hfe00;
			16'hd3b8: y = 16'hfe00;
			16'hd3b9: y = 16'hfe00;
			16'hd3ba: y = 16'hfe00;
			16'hd3bb: y = 16'hfe00;
			16'hd3bc: y = 16'hfe00;
			16'hd3bd: y = 16'hfe00;
			16'hd3be: y = 16'hfe00;
			16'hd3bf: y = 16'hfe00;
			16'hd3c0: y = 16'hfe00;
			16'hd3c1: y = 16'hfe00;
			16'hd3c2: y = 16'hfe00;
			16'hd3c3: y = 16'hfe00;
			16'hd3c4: y = 16'hfe00;
			16'hd3c5: y = 16'hfe00;
			16'hd3c6: y = 16'hfe00;
			16'hd3c7: y = 16'hfe00;
			16'hd3c8: y = 16'hfe00;
			16'hd3c9: y = 16'hfe00;
			16'hd3ca: y = 16'hfe00;
			16'hd3cb: y = 16'hfe00;
			16'hd3cc: y = 16'hfe00;
			16'hd3cd: y = 16'hfe00;
			16'hd3ce: y = 16'hfe00;
			16'hd3cf: y = 16'hfe00;
			16'hd3d0: y = 16'hfe00;
			16'hd3d1: y = 16'hfe00;
			16'hd3d2: y = 16'hfe00;
			16'hd3d3: y = 16'hfe00;
			16'hd3d4: y = 16'hfe00;
			16'hd3d5: y = 16'hfe00;
			16'hd3d6: y = 16'hfe00;
			16'hd3d7: y = 16'hfe00;
			16'hd3d8: y = 16'hfe00;
			16'hd3d9: y = 16'hfe00;
			16'hd3da: y = 16'hfe00;
			16'hd3db: y = 16'hfe00;
			16'hd3dc: y = 16'hfe00;
			16'hd3dd: y = 16'hfe00;
			16'hd3de: y = 16'hfe00;
			16'hd3df: y = 16'hfe00;
			16'hd3e0: y = 16'hfe00;
			16'hd3e1: y = 16'hfe00;
			16'hd3e2: y = 16'hfe00;
			16'hd3e3: y = 16'hfe00;
			16'hd3e4: y = 16'hfe00;
			16'hd3e5: y = 16'hfe00;
			16'hd3e6: y = 16'hfe00;
			16'hd3e7: y = 16'hfe00;
			16'hd3e8: y = 16'hfe00;
			16'hd3e9: y = 16'hfe00;
			16'hd3ea: y = 16'hfe00;
			16'hd3eb: y = 16'hfe00;
			16'hd3ec: y = 16'hfe00;
			16'hd3ed: y = 16'hfe00;
			16'hd3ee: y = 16'hfe00;
			16'hd3ef: y = 16'hfe00;
			16'hd3f0: y = 16'hfe00;
			16'hd3f1: y = 16'hfe00;
			16'hd3f2: y = 16'hfe00;
			16'hd3f3: y = 16'hfe00;
			16'hd3f4: y = 16'hfe00;
			16'hd3f5: y = 16'hfe00;
			16'hd3f6: y = 16'hfe00;
			16'hd3f7: y = 16'hfe00;
			16'hd3f8: y = 16'hfe00;
			16'hd3f9: y = 16'hfe00;
			16'hd3fa: y = 16'hfe00;
			16'hd3fb: y = 16'hfe00;
			16'hd3fc: y = 16'hfe00;
			16'hd3fd: y = 16'hfe00;
			16'hd3fe: y = 16'hfe00;
			16'hd3ff: y = 16'hfe00;
			16'hd400: y = 16'hfe00;
			16'hd401: y = 16'hfe00;
			16'hd402: y = 16'hfe00;
			16'hd403: y = 16'hfe00;
			16'hd404: y = 16'hfe00;
			16'hd405: y = 16'hfe00;
			16'hd406: y = 16'hfe00;
			16'hd407: y = 16'hfe00;
			16'hd408: y = 16'hfe00;
			16'hd409: y = 16'hfe00;
			16'hd40a: y = 16'hfe00;
			16'hd40b: y = 16'hfe00;
			16'hd40c: y = 16'hfe00;
			16'hd40d: y = 16'hfe00;
			16'hd40e: y = 16'hfe00;
			16'hd40f: y = 16'hfe00;
			16'hd410: y = 16'hfe00;
			16'hd411: y = 16'hfe00;
			16'hd412: y = 16'hfe00;
			16'hd413: y = 16'hfe00;
			16'hd414: y = 16'hfe00;
			16'hd415: y = 16'hfe00;
			16'hd416: y = 16'hfe00;
			16'hd417: y = 16'hfe00;
			16'hd418: y = 16'hfe00;
			16'hd419: y = 16'hfe00;
			16'hd41a: y = 16'hfe00;
			16'hd41b: y = 16'hfe00;
			16'hd41c: y = 16'hfe00;
			16'hd41d: y = 16'hfe00;
			16'hd41e: y = 16'hfe00;
			16'hd41f: y = 16'hfe00;
			16'hd420: y = 16'hfe00;
			16'hd421: y = 16'hfe00;
			16'hd422: y = 16'hfe00;
			16'hd423: y = 16'hfe00;
			16'hd424: y = 16'hfe00;
			16'hd425: y = 16'hfe00;
			16'hd426: y = 16'hfe00;
			16'hd427: y = 16'hfe00;
			16'hd428: y = 16'hfe00;
			16'hd429: y = 16'hfe00;
			16'hd42a: y = 16'hfe00;
			16'hd42b: y = 16'hfe00;
			16'hd42c: y = 16'hfe00;
			16'hd42d: y = 16'hfe00;
			16'hd42e: y = 16'hfe00;
			16'hd42f: y = 16'hfe00;
			16'hd430: y = 16'hfe00;
			16'hd431: y = 16'hfe00;
			16'hd432: y = 16'hfe00;
			16'hd433: y = 16'hfe00;
			16'hd434: y = 16'hfe00;
			16'hd435: y = 16'hfe00;
			16'hd436: y = 16'hfe00;
			16'hd437: y = 16'hfe00;
			16'hd438: y = 16'hfe00;
			16'hd439: y = 16'hfe00;
			16'hd43a: y = 16'hfe00;
			16'hd43b: y = 16'hfe00;
			16'hd43c: y = 16'hfe00;
			16'hd43d: y = 16'hfe00;
			16'hd43e: y = 16'hfe00;
			16'hd43f: y = 16'hfe00;
			16'hd440: y = 16'hfe00;
			16'hd441: y = 16'hfe00;
			16'hd442: y = 16'hfe00;
			16'hd443: y = 16'hfe00;
			16'hd444: y = 16'hfe00;
			16'hd445: y = 16'hfe00;
			16'hd446: y = 16'hfe00;
			16'hd447: y = 16'hfe00;
			16'hd448: y = 16'hfe00;
			16'hd449: y = 16'hfe00;
			16'hd44a: y = 16'hfe00;
			16'hd44b: y = 16'hfe00;
			16'hd44c: y = 16'hfe00;
			16'hd44d: y = 16'hfe00;
			16'hd44e: y = 16'hfe00;
			16'hd44f: y = 16'hfe00;
			16'hd450: y = 16'hfe00;
			16'hd451: y = 16'hfe00;
			16'hd452: y = 16'hfe00;
			16'hd453: y = 16'hfe00;
			16'hd454: y = 16'hfe00;
			16'hd455: y = 16'hfe00;
			16'hd456: y = 16'hfe00;
			16'hd457: y = 16'hfe00;
			16'hd458: y = 16'hfe00;
			16'hd459: y = 16'hfe00;
			16'hd45a: y = 16'hfe00;
			16'hd45b: y = 16'hfe00;
			16'hd45c: y = 16'hfe00;
			16'hd45d: y = 16'hfe00;
			16'hd45e: y = 16'hfe00;
			16'hd45f: y = 16'hfe00;
			16'hd460: y = 16'hfe00;
			16'hd461: y = 16'hfe00;
			16'hd462: y = 16'hfe00;
			16'hd463: y = 16'hfe00;
			16'hd464: y = 16'hfe00;
			16'hd465: y = 16'hfe00;
			16'hd466: y = 16'hfe00;
			16'hd467: y = 16'hfe00;
			16'hd468: y = 16'hfe00;
			16'hd469: y = 16'hfe00;
			16'hd46a: y = 16'hfe00;
			16'hd46b: y = 16'hfe00;
			16'hd46c: y = 16'hfe00;
			16'hd46d: y = 16'hfe00;
			16'hd46e: y = 16'hfe00;
			16'hd46f: y = 16'hfe00;
			16'hd470: y = 16'hfe00;
			16'hd471: y = 16'hfe00;
			16'hd472: y = 16'hfe00;
			16'hd473: y = 16'hfe00;
			16'hd474: y = 16'hfe00;
			16'hd475: y = 16'hfe00;
			16'hd476: y = 16'hfe00;
			16'hd477: y = 16'hfe00;
			16'hd478: y = 16'hfe00;
			16'hd479: y = 16'hfe00;
			16'hd47a: y = 16'hfe00;
			16'hd47b: y = 16'hfe00;
			16'hd47c: y = 16'hfe00;
			16'hd47d: y = 16'hfe00;
			16'hd47e: y = 16'hfe00;
			16'hd47f: y = 16'hfe00;
			16'hd480: y = 16'hfe00;
			16'hd481: y = 16'hfe00;
			16'hd482: y = 16'hfe00;
			16'hd483: y = 16'hfe00;
			16'hd484: y = 16'hfe00;
			16'hd485: y = 16'hfe00;
			16'hd486: y = 16'hfe00;
			16'hd487: y = 16'hfe00;
			16'hd488: y = 16'hfe00;
			16'hd489: y = 16'hfe00;
			16'hd48a: y = 16'hfe00;
			16'hd48b: y = 16'hfe00;
			16'hd48c: y = 16'hfe00;
			16'hd48d: y = 16'hfe00;
			16'hd48e: y = 16'hfe00;
			16'hd48f: y = 16'hfe00;
			16'hd490: y = 16'hfe00;
			16'hd491: y = 16'hfe00;
			16'hd492: y = 16'hfe00;
			16'hd493: y = 16'hfe00;
			16'hd494: y = 16'hfe00;
			16'hd495: y = 16'hfe00;
			16'hd496: y = 16'hfe00;
			16'hd497: y = 16'hfe00;
			16'hd498: y = 16'hfe00;
			16'hd499: y = 16'hfe00;
			16'hd49a: y = 16'hfe00;
			16'hd49b: y = 16'hfe00;
			16'hd49c: y = 16'hfe00;
			16'hd49d: y = 16'hfe00;
			16'hd49e: y = 16'hfe00;
			16'hd49f: y = 16'hfe00;
			16'hd4a0: y = 16'hfe00;
			16'hd4a1: y = 16'hfe00;
			16'hd4a2: y = 16'hfe00;
			16'hd4a3: y = 16'hfe00;
			16'hd4a4: y = 16'hfe00;
			16'hd4a5: y = 16'hfe00;
			16'hd4a6: y = 16'hfe00;
			16'hd4a7: y = 16'hfe00;
			16'hd4a8: y = 16'hfe00;
			16'hd4a9: y = 16'hfe00;
			16'hd4aa: y = 16'hfe00;
			16'hd4ab: y = 16'hfe00;
			16'hd4ac: y = 16'hfe00;
			16'hd4ad: y = 16'hfe00;
			16'hd4ae: y = 16'hfe00;
			16'hd4af: y = 16'hfe00;
			16'hd4b0: y = 16'hfe00;
			16'hd4b1: y = 16'hfe00;
			16'hd4b2: y = 16'hfe00;
			16'hd4b3: y = 16'hfe00;
			16'hd4b4: y = 16'hfe00;
			16'hd4b5: y = 16'hfe00;
			16'hd4b6: y = 16'hfe00;
			16'hd4b7: y = 16'hfe00;
			16'hd4b8: y = 16'hfe00;
			16'hd4b9: y = 16'hfe00;
			16'hd4ba: y = 16'hfe00;
			16'hd4bb: y = 16'hfe00;
			16'hd4bc: y = 16'hfe00;
			16'hd4bd: y = 16'hfe00;
			16'hd4be: y = 16'hfe00;
			16'hd4bf: y = 16'hfe00;
			16'hd4c0: y = 16'hfe00;
			16'hd4c1: y = 16'hfe00;
			16'hd4c2: y = 16'hfe00;
			16'hd4c3: y = 16'hfe00;
			16'hd4c4: y = 16'hfe00;
			16'hd4c5: y = 16'hfe00;
			16'hd4c6: y = 16'hfe00;
			16'hd4c7: y = 16'hfe00;
			16'hd4c8: y = 16'hfe00;
			16'hd4c9: y = 16'hfe00;
			16'hd4ca: y = 16'hfe00;
			16'hd4cb: y = 16'hfe00;
			16'hd4cc: y = 16'hfe00;
			16'hd4cd: y = 16'hfe00;
			16'hd4ce: y = 16'hfe00;
			16'hd4cf: y = 16'hfe00;
			16'hd4d0: y = 16'hfe00;
			16'hd4d1: y = 16'hfe00;
			16'hd4d2: y = 16'hfe00;
			16'hd4d3: y = 16'hfe00;
			16'hd4d4: y = 16'hfe00;
			16'hd4d5: y = 16'hfe00;
			16'hd4d6: y = 16'hfe00;
			16'hd4d7: y = 16'hfe00;
			16'hd4d8: y = 16'hfe00;
			16'hd4d9: y = 16'hfe00;
			16'hd4da: y = 16'hfe00;
			16'hd4db: y = 16'hfe00;
			16'hd4dc: y = 16'hfe00;
			16'hd4dd: y = 16'hfe00;
			16'hd4de: y = 16'hfe00;
			16'hd4df: y = 16'hfe00;
			16'hd4e0: y = 16'hfe00;
			16'hd4e1: y = 16'hfe00;
			16'hd4e2: y = 16'hfe00;
			16'hd4e3: y = 16'hfe00;
			16'hd4e4: y = 16'hfe00;
			16'hd4e5: y = 16'hfe00;
			16'hd4e6: y = 16'hfe00;
			16'hd4e7: y = 16'hfe00;
			16'hd4e8: y = 16'hfe00;
			16'hd4e9: y = 16'hfe00;
			16'hd4ea: y = 16'hfe00;
			16'hd4eb: y = 16'hfe00;
			16'hd4ec: y = 16'hfe00;
			16'hd4ed: y = 16'hfe00;
			16'hd4ee: y = 16'hfe00;
			16'hd4ef: y = 16'hfe00;
			16'hd4f0: y = 16'hfe00;
			16'hd4f1: y = 16'hfe00;
			16'hd4f2: y = 16'hfe00;
			16'hd4f3: y = 16'hfe00;
			16'hd4f4: y = 16'hfe00;
			16'hd4f5: y = 16'hfe00;
			16'hd4f6: y = 16'hfe00;
			16'hd4f7: y = 16'hfe00;
			16'hd4f8: y = 16'hfe00;
			16'hd4f9: y = 16'hfe00;
			16'hd4fa: y = 16'hfe00;
			16'hd4fb: y = 16'hfe00;
			16'hd4fc: y = 16'hfe00;
			16'hd4fd: y = 16'hfe00;
			16'hd4fe: y = 16'hfe00;
			16'hd4ff: y = 16'hfe00;
			16'hd500: y = 16'hfe00;
			16'hd501: y = 16'hfe00;
			16'hd502: y = 16'hfe00;
			16'hd503: y = 16'hfe00;
			16'hd504: y = 16'hfe00;
			16'hd505: y = 16'hfe00;
			16'hd506: y = 16'hfe00;
			16'hd507: y = 16'hfe00;
			16'hd508: y = 16'hfe00;
			16'hd509: y = 16'hfe00;
			16'hd50a: y = 16'hfe00;
			16'hd50b: y = 16'hfe00;
			16'hd50c: y = 16'hfe00;
			16'hd50d: y = 16'hfe00;
			16'hd50e: y = 16'hfe00;
			16'hd50f: y = 16'hfe00;
			16'hd510: y = 16'hfe00;
			16'hd511: y = 16'hfe00;
			16'hd512: y = 16'hfe00;
			16'hd513: y = 16'hfe00;
			16'hd514: y = 16'hfe00;
			16'hd515: y = 16'hfe00;
			16'hd516: y = 16'hfe00;
			16'hd517: y = 16'hfe00;
			16'hd518: y = 16'hfe00;
			16'hd519: y = 16'hfe00;
			16'hd51a: y = 16'hfe00;
			16'hd51b: y = 16'hfe00;
			16'hd51c: y = 16'hfe00;
			16'hd51d: y = 16'hfe00;
			16'hd51e: y = 16'hfe00;
			16'hd51f: y = 16'hfe00;
			16'hd520: y = 16'hfe00;
			16'hd521: y = 16'hfe00;
			16'hd522: y = 16'hfe00;
			16'hd523: y = 16'hfe00;
			16'hd524: y = 16'hfe00;
			16'hd525: y = 16'hfe00;
			16'hd526: y = 16'hfe00;
			16'hd527: y = 16'hfe00;
			16'hd528: y = 16'hfe00;
			16'hd529: y = 16'hfe00;
			16'hd52a: y = 16'hfe00;
			16'hd52b: y = 16'hfe00;
			16'hd52c: y = 16'hfe00;
			16'hd52d: y = 16'hfe00;
			16'hd52e: y = 16'hfe00;
			16'hd52f: y = 16'hfe00;
			16'hd530: y = 16'hfe00;
			16'hd531: y = 16'hfe00;
			16'hd532: y = 16'hfe00;
			16'hd533: y = 16'hfe00;
			16'hd534: y = 16'hfe00;
			16'hd535: y = 16'hfe00;
			16'hd536: y = 16'hfe00;
			16'hd537: y = 16'hfe00;
			16'hd538: y = 16'hfe00;
			16'hd539: y = 16'hfe00;
			16'hd53a: y = 16'hfe00;
			16'hd53b: y = 16'hfe00;
			16'hd53c: y = 16'hfe00;
			16'hd53d: y = 16'hfe00;
			16'hd53e: y = 16'hfe00;
			16'hd53f: y = 16'hfe00;
			16'hd540: y = 16'hfe00;
			16'hd541: y = 16'hfe00;
			16'hd542: y = 16'hfe00;
			16'hd543: y = 16'hfe00;
			16'hd544: y = 16'hfe00;
			16'hd545: y = 16'hfe00;
			16'hd546: y = 16'hfe00;
			16'hd547: y = 16'hfe00;
			16'hd548: y = 16'hfe00;
			16'hd549: y = 16'hfe00;
			16'hd54a: y = 16'hfe00;
			16'hd54b: y = 16'hfe00;
			16'hd54c: y = 16'hfe00;
			16'hd54d: y = 16'hfe00;
			16'hd54e: y = 16'hfe00;
			16'hd54f: y = 16'hfe00;
			16'hd550: y = 16'hfe00;
			16'hd551: y = 16'hfe00;
			16'hd552: y = 16'hfe00;
			16'hd553: y = 16'hfe00;
			16'hd554: y = 16'hfe00;
			16'hd555: y = 16'hfe00;
			16'hd556: y = 16'hfe00;
			16'hd557: y = 16'hfe00;
			16'hd558: y = 16'hfe00;
			16'hd559: y = 16'hfe00;
			16'hd55a: y = 16'hfe00;
			16'hd55b: y = 16'hfe00;
			16'hd55c: y = 16'hfe00;
			16'hd55d: y = 16'hfe00;
			16'hd55e: y = 16'hfe00;
			16'hd55f: y = 16'hfe00;
			16'hd560: y = 16'hfe00;
			16'hd561: y = 16'hfe00;
			16'hd562: y = 16'hfe00;
			16'hd563: y = 16'hfe00;
			16'hd564: y = 16'hfe00;
			16'hd565: y = 16'hfe00;
			16'hd566: y = 16'hfe00;
			16'hd567: y = 16'hfe00;
			16'hd568: y = 16'hfe00;
			16'hd569: y = 16'hfe00;
			16'hd56a: y = 16'hfe00;
			16'hd56b: y = 16'hfe00;
			16'hd56c: y = 16'hfe00;
			16'hd56d: y = 16'hfe00;
			16'hd56e: y = 16'hfe00;
			16'hd56f: y = 16'hfe00;
			16'hd570: y = 16'hfe00;
			16'hd571: y = 16'hfe00;
			16'hd572: y = 16'hfe00;
			16'hd573: y = 16'hfe00;
			16'hd574: y = 16'hfe00;
			16'hd575: y = 16'hfe00;
			16'hd576: y = 16'hfe00;
			16'hd577: y = 16'hfe00;
			16'hd578: y = 16'hfe00;
			16'hd579: y = 16'hfe00;
			16'hd57a: y = 16'hfe00;
			16'hd57b: y = 16'hfe00;
			16'hd57c: y = 16'hfe00;
			16'hd57d: y = 16'hfe00;
			16'hd57e: y = 16'hfe00;
			16'hd57f: y = 16'hfe00;
			16'hd580: y = 16'hfe00;
			16'hd581: y = 16'hfe00;
			16'hd582: y = 16'hfe00;
			16'hd583: y = 16'hfe00;
			16'hd584: y = 16'hfe00;
			16'hd585: y = 16'hfe00;
			16'hd586: y = 16'hfe00;
			16'hd587: y = 16'hfe00;
			16'hd588: y = 16'hfe00;
			16'hd589: y = 16'hfe00;
			16'hd58a: y = 16'hfe00;
			16'hd58b: y = 16'hfe00;
			16'hd58c: y = 16'hfe00;
			16'hd58d: y = 16'hfe00;
			16'hd58e: y = 16'hfe00;
			16'hd58f: y = 16'hfe00;
			16'hd590: y = 16'hfe00;
			16'hd591: y = 16'hfe00;
			16'hd592: y = 16'hfe00;
			16'hd593: y = 16'hfe00;
			16'hd594: y = 16'hfe00;
			16'hd595: y = 16'hfe00;
			16'hd596: y = 16'hfe00;
			16'hd597: y = 16'hfe00;
			16'hd598: y = 16'hfe00;
			16'hd599: y = 16'hfe00;
			16'hd59a: y = 16'hfe00;
			16'hd59b: y = 16'hfe00;
			16'hd59c: y = 16'hfe00;
			16'hd59d: y = 16'hfe00;
			16'hd59e: y = 16'hfe00;
			16'hd59f: y = 16'hfe00;
			16'hd5a0: y = 16'hfe00;
			16'hd5a1: y = 16'hfe00;
			16'hd5a2: y = 16'hfe00;
			16'hd5a3: y = 16'hfe00;
			16'hd5a4: y = 16'hfe00;
			16'hd5a5: y = 16'hfe00;
			16'hd5a6: y = 16'hfe00;
			16'hd5a7: y = 16'hfe00;
			16'hd5a8: y = 16'hfe00;
			16'hd5a9: y = 16'hfe00;
			16'hd5aa: y = 16'hfe00;
			16'hd5ab: y = 16'hfe00;
			16'hd5ac: y = 16'hfe00;
			16'hd5ad: y = 16'hfe00;
			16'hd5ae: y = 16'hfe00;
			16'hd5af: y = 16'hfe00;
			16'hd5b0: y = 16'hfe00;
			16'hd5b1: y = 16'hfe00;
			16'hd5b2: y = 16'hfe00;
			16'hd5b3: y = 16'hfe00;
			16'hd5b4: y = 16'hfe00;
			16'hd5b5: y = 16'hfe00;
			16'hd5b6: y = 16'hfe00;
			16'hd5b7: y = 16'hfe00;
			16'hd5b8: y = 16'hfe00;
			16'hd5b9: y = 16'hfe00;
			16'hd5ba: y = 16'hfe00;
			16'hd5bb: y = 16'hfe00;
			16'hd5bc: y = 16'hfe00;
			16'hd5bd: y = 16'hfe00;
			16'hd5be: y = 16'hfe00;
			16'hd5bf: y = 16'hfe00;
			16'hd5c0: y = 16'hfe00;
			16'hd5c1: y = 16'hfe00;
			16'hd5c2: y = 16'hfe00;
			16'hd5c3: y = 16'hfe00;
			16'hd5c4: y = 16'hfe00;
			16'hd5c5: y = 16'hfe00;
			16'hd5c6: y = 16'hfe00;
			16'hd5c7: y = 16'hfe00;
			16'hd5c8: y = 16'hfe00;
			16'hd5c9: y = 16'hfe00;
			16'hd5ca: y = 16'hfe00;
			16'hd5cb: y = 16'hfe00;
			16'hd5cc: y = 16'hfe00;
			16'hd5cd: y = 16'hfe00;
			16'hd5ce: y = 16'hfe00;
			16'hd5cf: y = 16'hfe00;
			16'hd5d0: y = 16'hfe00;
			16'hd5d1: y = 16'hfe00;
			16'hd5d2: y = 16'hfe00;
			16'hd5d3: y = 16'hfe00;
			16'hd5d4: y = 16'hfe00;
			16'hd5d5: y = 16'hfe00;
			16'hd5d6: y = 16'hfe00;
			16'hd5d7: y = 16'hfe00;
			16'hd5d8: y = 16'hfe00;
			16'hd5d9: y = 16'hfe00;
			16'hd5da: y = 16'hfe00;
			16'hd5db: y = 16'hfe00;
			16'hd5dc: y = 16'hfe00;
			16'hd5dd: y = 16'hfe00;
			16'hd5de: y = 16'hfe00;
			16'hd5df: y = 16'hfe00;
			16'hd5e0: y = 16'hfe00;
			16'hd5e1: y = 16'hfe00;
			16'hd5e2: y = 16'hfe00;
			16'hd5e3: y = 16'hfe00;
			16'hd5e4: y = 16'hfe00;
			16'hd5e5: y = 16'hfe00;
			16'hd5e6: y = 16'hfe00;
			16'hd5e7: y = 16'hfe00;
			16'hd5e8: y = 16'hfe00;
			16'hd5e9: y = 16'hfe00;
			16'hd5ea: y = 16'hfe00;
			16'hd5eb: y = 16'hfe00;
			16'hd5ec: y = 16'hfe00;
			16'hd5ed: y = 16'hfe00;
			16'hd5ee: y = 16'hfe00;
			16'hd5ef: y = 16'hfe00;
			16'hd5f0: y = 16'hfe00;
			16'hd5f1: y = 16'hfe00;
			16'hd5f2: y = 16'hfe00;
			16'hd5f3: y = 16'hfe00;
			16'hd5f4: y = 16'hfe00;
			16'hd5f5: y = 16'hfe00;
			16'hd5f6: y = 16'hfe00;
			16'hd5f7: y = 16'hfe00;
			16'hd5f8: y = 16'hfe00;
			16'hd5f9: y = 16'hfe00;
			16'hd5fa: y = 16'hfe00;
			16'hd5fb: y = 16'hfe00;
			16'hd5fc: y = 16'hfe00;
			16'hd5fd: y = 16'hfe00;
			16'hd5fe: y = 16'hfe00;
			16'hd5ff: y = 16'hfe00;
			16'hd600: y = 16'hfe00;
			16'hd601: y = 16'hfe00;
			16'hd602: y = 16'hfe00;
			16'hd603: y = 16'hfe00;
			16'hd604: y = 16'hfe00;
			16'hd605: y = 16'hfe00;
			16'hd606: y = 16'hfe00;
			16'hd607: y = 16'hfe00;
			16'hd608: y = 16'hfe00;
			16'hd609: y = 16'hfe00;
			16'hd60a: y = 16'hfe00;
			16'hd60b: y = 16'hfe00;
			16'hd60c: y = 16'hfe00;
			16'hd60d: y = 16'hfe00;
			16'hd60e: y = 16'hfe00;
			16'hd60f: y = 16'hfe00;
			16'hd610: y = 16'hfe00;
			16'hd611: y = 16'hfe00;
			16'hd612: y = 16'hfe00;
			16'hd613: y = 16'hfe00;
			16'hd614: y = 16'hfe00;
			16'hd615: y = 16'hfe00;
			16'hd616: y = 16'hfe00;
			16'hd617: y = 16'hfe00;
			16'hd618: y = 16'hfe00;
			16'hd619: y = 16'hfe00;
			16'hd61a: y = 16'hfe00;
			16'hd61b: y = 16'hfe00;
			16'hd61c: y = 16'hfe00;
			16'hd61d: y = 16'hfe00;
			16'hd61e: y = 16'hfe00;
			16'hd61f: y = 16'hfe00;
			16'hd620: y = 16'hfe00;
			16'hd621: y = 16'hfe00;
			16'hd622: y = 16'hfe00;
			16'hd623: y = 16'hfe00;
			16'hd624: y = 16'hfe00;
			16'hd625: y = 16'hfe00;
			16'hd626: y = 16'hfe00;
			16'hd627: y = 16'hfe00;
			16'hd628: y = 16'hfe00;
			16'hd629: y = 16'hfe00;
			16'hd62a: y = 16'hfe00;
			16'hd62b: y = 16'hfe00;
			16'hd62c: y = 16'hfe00;
			16'hd62d: y = 16'hfe00;
			16'hd62e: y = 16'hfe00;
			16'hd62f: y = 16'hfe00;
			16'hd630: y = 16'hfe00;
			16'hd631: y = 16'hfe00;
			16'hd632: y = 16'hfe00;
			16'hd633: y = 16'hfe00;
			16'hd634: y = 16'hfe00;
			16'hd635: y = 16'hfe00;
			16'hd636: y = 16'hfe00;
			16'hd637: y = 16'hfe00;
			16'hd638: y = 16'hfe00;
			16'hd639: y = 16'hfe00;
			16'hd63a: y = 16'hfe00;
			16'hd63b: y = 16'hfe00;
			16'hd63c: y = 16'hfe00;
			16'hd63d: y = 16'hfe00;
			16'hd63e: y = 16'hfe00;
			16'hd63f: y = 16'hfe00;
			16'hd640: y = 16'hfe00;
			16'hd641: y = 16'hfe00;
			16'hd642: y = 16'hfe00;
			16'hd643: y = 16'hfe00;
			16'hd644: y = 16'hfe00;
			16'hd645: y = 16'hfe00;
			16'hd646: y = 16'hfe00;
			16'hd647: y = 16'hfe00;
			16'hd648: y = 16'hfe00;
			16'hd649: y = 16'hfe00;
			16'hd64a: y = 16'hfe00;
			16'hd64b: y = 16'hfe00;
			16'hd64c: y = 16'hfe00;
			16'hd64d: y = 16'hfe00;
			16'hd64e: y = 16'hfe00;
			16'hd64f: y = 16'hfe00;
			16'hd650: y = 16'hfe00;
			16'hd651: y = 16'hfe00;
			16'hd652: y = 16'hfe00;
			16'hd653: y = 16'hfe00;
			16'hd654: y = 16'hfe00;
			16'hd655: y = 16'hfe00;
			16'hd656: y = 16'hfe00;
			16'hd657: y = 16'hfe00;
			16'hd658: y = 16'hfe00;
			16'hd659: y = 16'hfe00;
			16'hd65a: y = 16'hfe00;
			16'hd65b: y = 16'hfe00;
			16'hd65c: y = 16'hfe00;
			16'hd65d: y = 16'hfe00;
			16'hd65e: y = 16'hfe00;
			16'hd65f: y = 16'hfe00;
			16'hd660: y = 16'hfe00;
			16'hd661: y = 16'hfe00;
			16'hd662: y = 16'hfe00;
			16'hd663: y = 16'hfe00;
			16'hd664: y = 16'hfe00;
			16'hd665: y = 16'hfe00;
			16'hd666: y = 16'hfe00;
			16'hd667: y = 16'hfe00;
			16'hd668: y = 16'hfe00;
			16'hd669: y = 16'hfe00;
			16'hd66a: y = 16'hfe00;
			16'hd66b: y = 16'hfe00;
			16'hd66c: y = 16'hfe00;
			16'hd66d: y = 16'hfe00;
			16'hd66e: y = 16'hfe00;
			16'hd66f: y = 16'hfe00;
			16'hd670: y = 16'hfe00;
			16'hd671: y = 16'hfe00;
			16'hd672: y = 16'hfe00;
			16'hd673: y = 16'hfe00;
			16'hd674: y = 16'hfe00;
			16'hd675: y = 16'hfe00;
			16'hd676: y = 16'hfe00;
			16'hd677: y = 16'hfe00;
			16'hd678: y = 16'hfe00;
			16'hd679: y = 16'hfe00;
			16'hd67a: y = 16'hfe00;
			16'hd67b: y = 16'hfe00;
			16'hd67c: y = 16'hfe00;
			16'hd67d: y = 16'hfe00;
			16'hd67e: y = 16'hfe00;
			16'hd67f: y = 16'hfe00;
			16'hd680: y = 16'hfe00;
			16'hd681: y = 16'hfe00;
			16'hd682: y = 16'hfe00;
			16'hd683: y = 16'hfe00;
			16'hd684: y = 16'hfe00;
			16'hd685: y = 16'hfe00;
			16'hd686: y = 16'hfe00;
			16'hd687: y = 16'hfe00;
			16'hd688: y = 16'hfe00;
			16'hd689: y = 16'hfe00;
			16'hd68a: y = 16'hfe00;
			16'hd68b: y = 16'hfe00;
			16'hd68c: y = 16'hfe00;
			16'hd68d: y = 16'hfe00;
			16'hd68e: y = 16'hfe00;
			16'hd68f: y = 16'hfe00;
			16'hd690: y = 16'hfe00;
			16'hd691: y = 16'hfe00;
			16'hd692: y = 16'hfe00;
			16'hd693: y = 16'hfe00;
			16'hd694: y = 16'hfe00;
			16'hd695: y = 16'hfe00;
			16'hd696: y = 16'hfe00;
			16'hd697: y = 16'hfe00;
			16'hd698: y = 16'hfe00;
			16'hd699: y = 16'hfe00;
			16'hd69a: y = 16'hfe00;
			16'hd69b: y = 16'hfe00;
			16'hd69c: y = 16'hfe00;
			16'hd69d: y = 16'hfe00;
			16'hd69e: y = 16'hfe00;
			16'hd69f: y = 16'hfe00;
			16'hd6a0: y = 16'hfe00;
			16'hd6a1: y = 16'hfe00;
			16'hd6a2: y = 16'hfe00;
			16'hd6a3: y = 16'hfe00;
			16'hd6a4: y = 16'hfe00;
			16'hd6a5: y = 16'hfe00;
			16'hd6a6: y = 16'hfe00;
			16'hd6a7: y = 16'hfe00;
			16'hd6a8: y = 16'hfe00;
			16'hd6a9: y = 16'hfe00;
			16'hd6aa: y = 16'hfe00;
			16'hd6ab: y = 16'hfe00;
			16'hd6ac: y = 16'hfe00;
			16'hd6ad: y = 16'hfe00;
			16'hd6ae: y = 16'hfe00;
			16'hd6af: y = 16'hfe00;
			16'hd6b0: y = 16'hfe00;
			16'hd6b1: y = 16'hfe00;
			16'hd6b2: y = 16'hfe00;
			16'hd6b3: y = 16'hfe00;
			16'hd6b4: y = 16'hfe00;
			16'hd6b5: y = 16'hfe00;
			16'hd6b6: y = 16'hfe00;
			16'hd6b7: y = 16'hfe00;
			16'hd6b8: y = 16'hfe00;
			16'hd6b9: y = 16'hfe00;
			16'hd6ba: y = 16'hfe00;
			16'hd6bb: y = 16'hfe00;
			16'hd6bc: y = 16'hfe00;
			16'hd6bd: y = 16'hfe00;
			16'hd6be: y = 16'hfe00;
			16'hd6bf: y = 16'hfe00;
			16'hd6c0: y = 16'hfe00;
			16'hd6c1: y = 16'hfe00;
			16'hd6c2: y = 16'hfe00;
			16'hd6c3: y = 16'hfe00;
			16'hd6c4: y = 16'hfe00;
			16'hd6c5: y = 16'hfe00;
			16'hd6c6: y = 16'hfe00;
			16'hd6c7: y = 16'hfe00;
			16'hd6c8: y = 16'hfe00;
			16'hd6c9: y = 16'hfe00;
			16'hd6ca: y = 16'hfe00;
			16'hd6cb: y = 16'hfe00;
			16'hd6cc: y = 16'hfe00;
			16'hd6cd: y = 16'hfe00;
			16'hd6ce: y = 16'hfe00;
			16'hd6cf: y = 16'hfe00;
			16'hd6d0: y = 16'hfe00;
			16'hd6d1: y = 16'hfe00;
			16'hd6d2: y = 16'hfe00;
			16'hd6d3: y = 16'hfe00;
			16'hd6d4: y = 16'hfe00;
			16'hd6d5: y = 16'hfe00;
			16'hd6d6: y = 16'hfe00;
			16'hd6d7: y = 16'hfe00;
			16'hd6d8: y = 16'hfe00;
			16'hd6d9: y = 16'hfe00;
			16'hd6da: y = 16'hfe00;
			16'hd6db: y = 16'hfe00;
			16'hd6dc: y = 16'hfe00;
			16'hd6dd: y = 16'hfe00;
			16'hd6de: y = 16'hfe00;
			16'hd6df: y = 16'hfe00;
			16'hd6e0: y = 16'hfe00;
			16'hd6e1: y = 16'hfe00;
			16'hd6e2: y = 16'hfe00;
			16'hd6e3: y = 16'hfe00;
			16'hd6e4: y = 16'hfe00;
			16'hd6e5: y = 16'hfe00;
			16'hd6e6: y = 16'hfe00;
			16'hd6e7: y = 16'hfe00;
			16'hd6e8: y = 16'hfe00;
			16'hd6e9: y = 16'hfe00;
			16'hd6ea: y = 16'hfe00;
			16'hd6eb: y = 16'hfe00;
			16'hd6ec: y = 16'hfe00;
			16'hd6ed: y = 16'hfe00;
			16'hd6ee: y = 16'hfe00;
			16'hd6ef: y = 16'hfe00;
			16'hd6f0: y = 16'hfe00;
			16'hd6f1: y = 16'hfe00;
			16'hd6f2: y = 16'hfe00;
			16'hd6f3: y = 16'hfe00;
			16'hd6f4: y = 16'hfe00;
			16'hd6f5: y = 16'hfe00;
			16'hd6f6: y = 16'hfe00;
			16'hd6f7: y = 16'hfe00;
			16'hd6f8: y = 16'hfe00;
			16'hd6f9: y = 16'hfe00;
			16'hd6fa: y = 16'hfe00;
			16'hd6fb: y = 16'hfe00;
			16'hd6fc: y = 16'hfe00;
			16'hd6fd: y = 16'hfe00;
			16'hd6fe: y = 16'hfe00;
			16'hd6ff: y = 16'hfe00;
			16'hd700: y = 16'hfe00;
			16'hd701: y = 16'hfe00;
			16'hd702: y = 16'hfe00;
			16'hd703: y = 16'hfe00;
			16'hd704: y = 16'hfe00;
			16'hd705: y = 16'hfe00;
			16'hd706: y = 16'hfe00;
			16'hd707: y = 16'hfe00;
			16'hd708: y = 16'hfe00;
			16'hd709: y = 16'hfe00;
			16'hd70a: y = 16'hfe00;
			16'hd70b: y = 16'hfe00;
			16'hd70c: y = 16'hfe00;
			16'hd70d: y = 16'hfe00;
			16'hd70e: y = 16'hfe00;
			16'hd70f: y = 16'hfe00;
			16'hd710: y = 16'hfe00;
			16'hd711: y = 16'hfe00;
			16'hd712: y = 16'hfe00;
			16'hd713: y = 16'hfe00;
			16'hd714: y = 16'hfe00;
			16'hd715: y = 16'hfe00;
			16'hd716: y = 16'hfe00;
			16'hd717: y = 16'hfe00;
			16'hd718: y = 16'hfe00;
			16'hd719: y = 16'hfe00;
			16'hd71a: y = 16'hfe00;
			16'hd71b: y = 16'hfe00;
			16'hd71c: y = 16'hfe00;
			16'hd71d: y = 16'hfe00;
			16'hd71e: y = 16'hfe00;
			16'hd71f: y = 16'hfe00;
			16'hd720: y = 16'hfe00;
			16'hd721: y = 16'hfe00;
			16'hd722: y = 16'hfe00;
			16'hd723: y = 16'hfe00;
			16'hd724: y = 16'hfe00;
			16'hd725: y = 16'hfe00;
			16'hd726: y = 16'hfe00;
			16'hd727: y = 16'hfe00;
			16'hd728: y = 16'hfe00;
			16'hd729: y = 16'hfe00;
			16'hd72a: y = 16'hfe00;
			16'hd72b: y = 16'hfe00;
			16'hd72c: y = 16'hfe00;
			16'hd72d: y = 16'hfe00;
			16'hd72e: y = 16'hfe00;
			16'hd72f: y = 16'hfe00;
			16'hd730: y = 16'hfe00;
			16'hd731: y = 16'hfe00;
			16'hd732: y = 16'hfe00;
			16'hd733: y = 16'hfe00;
			16'hd734: y = 16'hfe00;
			16'hd735: y = 16'hfe00;
			16'hd736: y = 16'hfe00;
			16'hd737: y = 16'hfe00;
			16'hd738: y = 16'hfe00;
			16'hd739: y = 16'hfe00;
			16'hd73a: y = 16'hfe00;
			16'hd73b: y = 16'hfe00;
			16'hd73c: y = 16'hfe00;
			16'hd73d: y = 16'hfe00;
			16'hd73e: y = 16'hfe00;
			16'hd73f: y = 16'hfe00;
			16'hd740: y = 16'hfe00;
			16'hd741: y = 16'hfe00;
			16'hd742: y = 16'hfe00;
			16'hd743: y = 16'hfe00;
			16'hd744: y = 16'hfe00;
			16'hd745: y = 16'hfe00;
			16'hd746: y = 16'hfe00;
			16'hd747: y = 16'hfe00;
			16'hd748: y = 16'hfe00;
			16'hd749: y = 16'hfe00;
			16'hd74a: y = 16'hfe00;
			16'hd74b: y = 16'hfe00;
			16'hd74c: y = 16'hfe00;
			16'hd74d: y = 16'hfe00;
			16'hd74e: y = 16'hfe00;
			16'hd74f: y = 16'hfe00;
			16'hd750: y = 16'hfe00;
			16'hd751: y = 16'hfe00;
			16'hd752: y = 16'hfe00;
			16'hd753: y = 16'hfe00;
			16'hd754: y = 16'hfe00;
			16'hd755: y = 16'hfe00;
			16'hd756: y = 16'hfe00;
			16'hd757: y = 16'hfe00;
			16'hd758: y = 16'hfe00;
			16'hd759: y = 16'hfe00;
			16'hd75a: y = 16'hfe00;
			16'hd75b: y = 16'hfe00;
			16'hd75c: y = 16'hfe00;
			16'hd75d: y = 16'hfe00;
			16'hd75e: y = 16'hfe00;
			16'hd75f: y = 16'hfe00;
			16'hd760: y = 16'hfe00;
			16'hd761: y = 16'hfe00;
			16'hd762: y = 16'hfe00;
			16'hd763: y = 16'hfe00;
			16'hd764: y = 16'hfe00;
			16'hd765: y = 16'hfe00;
			16'hd766: y = 16'hfe00;
			16'hd767: y = 16'hfe00;
			16'hd768: y = 16'hfe00;
			16'hd769: y = 16'hfe00;
			16'hd76a: y = 16'hfe00;
			16'hd76b: y = 16'hfe00;
			16'hd76c: y = 16'hfe00;
			16'hd76d: y = 16'hfe00;
			16'hd76e: y = 16'hfe00;
			16'hd76f: y = 16'hfe00;
			16'hd770: y = 16'hfe00;
			16'hd771: y = 16'hfe00;
			16'hd772: y = 16'hfe00;
			16'hd773: y = 16'hfe00;
			16'hd774: y = 16'hfe00;
			16'hd775: y = 16'hfe00;
			16'hd776: y = 16'hfe00;
			16'hd777: y = 16'hfe00;
			16'hd778: y = 16'hfe00;
			16'hd779: y = 16'hfe00;
			16'hd77a: y = 16'hfe00;
			16'hd77b: y = 16'hfe00;
			16'hd77c: y = 16'hfe00;
			16'hd77d: y = 16'hfe00;
			16'hd77e: y = 16'hfe00;
			16'hd77f: y = 16'hfe00;
			16'hd780: y = 16'hfe00;
			16'hd781: y = 16'hfe00;
			16'hd782: y = 16'hfe00;
			16'hd783: y = 16'hfe00;
			16'hd784: y = 16'hfe00;
			16'hd785: y = 16'hfe00;
			16'hd786: y = 16'hfe00;
			16'hd787: y = 16'hfe00;
			16'hd788: y = 16'hfe00;
			16'hd789: y = 16'hfe00;
			16'hd78a: y = 16'hfe00;
			16'hd78b: y = 16'hfe00;
			16'hd78c: y = 16'hfe00;
			16'hd78d: y = 16'hfe00;
			16'hd78e: y = 16'hfe00;
			16'hd78f: y = 16'hfe00;
			16'hd790: y = 16'hfe00;
			16'hd791: y = 16'hfe00;
			16'hd792: y = 16'hfe00;
			16'hd793: y = 16'hfe00;
			16'hd794: y = 16'hfe00;
			16'hd795: y = 16'hfe00;
			16'hd796: y = 16'hfe00;
			16'hd797: y = 16'hfe00;
			16'hd798: y = 16'hfe00;
			16'hd799: y = 16'hfe00;
			16'hd79a: y = 16'hfe00;
			16'hd79b: y = 16'hfe00;
			16'hd79c: y = 16'hfe00;
			16'hd79d: y = 16'hfe00;
			16'hd79e: y = 16'hfe00;
			16'hd79f: y = 16'hfe00;
			16'hd7a0: y = 16'hfe00;
			16'hd7a1: y = 16'hfe00;
			16'hd7a2: y = 16'hfe00;
			16'hd7a3: y = 16'hfe00;
			16'hd7a4: y = 16'hfe00;
			16'hd7a5: y = 16'hfe00;
			16'hd7a6: y = 16'hfe00;
			16'hd7a7: y = 16'hfe00;
			16'hd7a8: y = 16'hfe00;
			16'hd7a9: y = 16'hfe00;
			16'hd7aa: y = 16'hfe00;
			16'hd7ab: y = 16'hfe00;
			16'hd7ac: y = 16'hfe00;
			16'hd7ad: y = 16'hfe00;
			16'hd7ae: y = 16'hfe00;
			16'hd7af: y = 16'hfe00;
			16'hd7b0: y = 16'hfe00;
			16'hd7b1: y = 16'hfe00;
			16'hd7b2: y = 16'hfe00;
			16'hd7b3: y = 16'hfe00;
			16'hd7b4: y = 16'hfe00;
			16'hd7b5: y = 16'hfe00;
			16'hd7b6: y = 16'hfe00;
			16'hd7b7: y = 16'hfe00;
			16'hd7b8: y = 16'hfe00;
			16'hd7b9: y = 16'hfe00;
			16'hd7ba: y = 16'hfe00;
			16'hd7bb: y = 16'hfe00;
			16'hd7bc: y = 16'hfe00;
			16'hd7bd: y = 16'hfe00;
			16'hd7be: y = 16'hfe00;
			16'hd7bf: y = 16'hfe00;
			16'hd7c0: y = 16'hfe00;
			16'hd7c1: y = 16'hfe00;
			16'hd7c2: y = 16'hfe00;
			16'hd7c3: y = 16'hfe00;
			16'hd7c4: y = 16'hfe00;
			16'hd7c5: y = 16'hfe00;
			16'hd7c6: y = 16'hfe00;
			16'hd7c7: y = 16'hfe00;
			16'hd7c8: y = 16'hfe00;
			16'hd7c9: y = 16'hfe00;
			16'hd7ca: y = 16'hfe00;
			16'hd7cb: y = 16'hfe00;
			16'hd7cc: y = 16'hfe00;
			16'hd7cd: y = 16'hfe00;
			16'hd7ce: y = 16'hfe00;
			16'hd7cf: y = 16'hfe00;
			16'hd7d0: y = 16'hfe00;
			16'hd7d1: y = 16'hfe00;
			16'hd7d2: y = 16'hfe00;
			16'hd7d3: y = 16'hfe00;
			16'hd7d4: y = 16'hfe00;
			16'hd7d5: y = 16'hfe00;
			16'hd7d6: y = 16'hfe00;
			16'hd7d7: y = 16'hfe00;
			16'hd7d8: y = 16'hfe00;
			16'hd7d9: y = 16'hfe00;
			16'hd7da: y = 16'hfe00;
			16'hd7db: y = 16'hfe00;
			16'hd7dc: y = 16'hfe00;
			16'hd7dd: y = 16'hfe00;
			16'hd7de: y = 16'hfe00;
			16'hd7df: y = 16'hfe00;
			16'hd7e0: y = 16'hfe00;
			16'hd7e1: y = 16'hfe00;
			16'hd7e2: y = 16'hfe00;
			16'hd7e3: y = 16'hfe00;
			16'hd7e4: y = 16'hfe00;
			16'hd7e5: y = 16'hfe00;
			16'hd7e6: y = 16'hfe00;
			16'hd7e7: y = 16'hfe00;
			16'hd7e8: y = 16'hfe00;
			16'hd7e9: y = 16'hfe00;
			16'hd7ea: y = 16'hfe00;
			16'hd7eb: y = 16'hfe00;
			16'hd7ec: y = 16'hfe00;
			16'hd7ed: y = 16'hfe00;
			16'hd7ee: y = 16'hfe00;
			16'hd7ef: y = 16'hfe00;
			16'hd7f0: y = 16'hfe00;
			16'hd7f1: y = 16'hfe00;
			16'hd7f2: y = 16'hfe00;
			16'hd7f3: y = 16'hfe00;
			16'hd7f4: y = 16'hfe00;
			16'hd7f5: y = 16'hfe00;
			16'hd7f6: y = 16'hfe00;
			16'hd7f7: y = 16'hfe00;
			16'hd7f8: y = 16'hfe00;
			16'hd7f9: y = 16'hfe00;
			16'hd7fa: y = 16'hfe00;
			16'hd7fb: y = 16'hfe00;
			16'hd7fc: y = 16'hfe00;
			16'hd7fd: y = 16'hfe00;
			16'hd7fe: y = 16'hfe00;
			16'hd7ff: y = 16'hfe00;
			16'hd800: y = 16'hfe00;
			16'hd801: y = 16'hfe00;
			16'hd802: y = 16'hfe00;
			16'hd803: y = 16'hfe00;
			16'hd804: y = 16'hfe00;
			16'hd805: y = 16'hfe00;
			16'hd806: y = 16'hfe00;
			16'hd807: y = 16'hfe00;
			16'hd808: y = 16'hfe00;
			16'hd809: y = 16'hfe00;
			16'hd80a: y = 16'hfe00;
			16'hd80b: y = 16'hfe00;
			16'hd80c: y = 16'hfe00;
			16'hd80d: y = 16'hfe00;
			16'hd80e: y = 16'hfe00;
			16'hd80f: y = 16'hfe00;
			16'hd810: y = 16'hfe00;
			16'hd811: y = 16'hfe00;
			16'hd812: y = 16'hfe00;
			16'hd813: y = 16'hfe00;
			16'hd814: y = 16'hfe00;
			16'hd815: y = 16'hfe00;
			16'hd816: y = 16'hfe00;
			16'hd817: y = 16'hfe00;
			16'hd818: y = 16'hfe00;
			16'hd819: y = 16'hfe00;
			16'hd81a: y = 16'hfe00;
			16'hd81b: y = 16'hfe00;
			16'hd81c: y = 16'hfe00;
			16'hd81d: y = 16'hfe00;
			16'hd81e: y = 16'hfe00;
			16'hd81f: y = 16'hfe00;
			16'hd820: y = 16'hfe00;
			16'hd821: y = 16'hfe00;
			16'hd822: y = 16'hfe00;
			16'hd823: y = 16'hfe00;
			16'hd824: y = 16'hfe00;
			16'hd825: y = 16'hfe00;
			16'hd826: y = 16'hfe00;
			16'hd827: y = 16'hfe00;
			16'hd828: y = 16'hfe00;
			16'hd829: y = 16'hfe00;
			16'hd82a: y = 16'hfe00;
			16'hd82b: y = 16'hfe00;
			16'hd82c: y = 16'hfe00;
			16'hd82d: y = 16'hfe00;
			16'hd82e: y = 16'hfe00;
			16'hd82f: y = 16'hfe00;
			16'hd830: y = 16'hfe00;
			16'hd831: y = 16'hfe00;
			16'hd832: y = 16'hfe00;
			16'hd833: y = 16'hfe00;
			16'hd834: y = 16'hfe00;
			16'hd835: y = 16'hfe00;
			16'hd836: y = 16'hfe00;
			16'hd837: y = 16'hfe00;
			16'hd838: y = 16'hfe00;
			16'hd839: y = 16'hfe00;
			16'hd83a: y = 16'hfe00;
			16'hd83b: y = 16'hfe00;
			16'hd83c: y = 16'hfe00;
			16'hd83d: y = 16'hfe00;
			16'hd83e: y = 16'hfe00;
			16'hd83f: y = 16'hfe00;
			16'hd840: y = 16'hfe00;
			16'hd841: y = 16'hfe00;
			16'hd842: y = 16'hfe00;
			16'hd843: y = 16'hfe00;
			16'hd844: y = 16'hfe00;
			16'hd845: y = 16'hfe00;
			16'hd846: y = 16'hfe00;
			16'hd847: y = 16'hfe00;
			16'hd848: y = 16'hfe00;
			16'hd849: y = 16'hfe00;
			16'hd84a: y = 16'hfe00;
			16'hd84b: y = 16'hfe00;
			16'hd84c: y = 16'hfe00;
			16'hd84d: y = 16'hfe00;
			16'hd84e: y = 16'hfe00;
			16'hd84f: y = 16'hfe00;
			16'hd850: y = 16'hfe00;
			16'hd851: y = 16'hfe00;
			16'hd852: y = 16'hfe00;
			16'hd853: y = 16'hfe00;
			16'hd854: y = 16'hfe00;
			16'hd855: y = 16'hfe00;
			16'hd856: y = 16'hfe00;
			16'hd857: y = 16'hfe00;
			16'hd858: y = 16'hfe00;
			16'hd859: y = 16'hfe00;
			16'hd85a: y = 16'hfe00;
			16'hd85b: y = 16'hfe00;
			16'hd85c: y = 16'hfe00;
			16'hd85d: y = 16'hfe00;
			16'hd85e: y = 16'hfe00;
			16'hd85f: y = 16'hfe00;
			16'hd860: y = 16'hfe00;
			16'hd861: y = 16'hfe00;
			16'hd862: y = 16'hfe00;
			16'hd863: y = 16'hfe00;
			16'hd864: y = 16'hfe00;
			16'hd865: y = 16'hfe00;
			16'hd866: y = 16'hfe00;
			16'hd867: y = 16'hfe00;
			16'hd868: y = 16'hfe00;
			16'hd869: y = 16'hfe00;
			16'hd86a: y = 16'hfe00;
			16'hd86b: y = 16'hfe00;
			16'hd86c: y = 16'hfe00;
			16'hd86d: y = 16'hfe00;
			16'hd86e: y = 16'hfe00;
			16'hd86f: y = 16'hfe00;
			16'hd870: y = 16'hfe00;
			16'hd871: y = 16'hfe00;
			16'hd872: y = 16'hfe00;
			16'hd873: y = 16'hfe00;
			16'hd874: y = 16'hfe00;
			16'hd875: y = 16'hfe00;
			16'hd876: y = 16'hfe00;
			16'hd877: y = 16'hfe00;
			16'hd878: y = 16'hfe00;
			16'hd879: y = 16'hfe00;
			16'hd87a: y = 16'hfe00;
			16'hd87b: y = 16'hfe00;
			16'hd87c: y = 16'hfe00;
			16'hd87d: y = 16'hfe00;
			16'hd87e: y = 16'hfe00;
			16'hd87f: y = 16'hfe00;
			16'hd880: y = 16'hfe00;
			16'hd881: y = 16'hfe00;
			16'hd882: y = 16'hfe00;
			16'hd883: y = 16'hfe00;
			16'hd884: y = 16'hfe00;
			16'hd885: y = 16'hfe00;
			16'hd886: y = 16'hfe00;
			16'hd887: y = 16'hfe00;
			16'hd888: y = 16'hfe00;
			16'hd889: y = 16'hfe00;
			16'hd88a: y = 16'hfe00;
			16'hd88b: y = 16'hfe00;
			16'hd88c: y = 16'hfe00;
			16'hd88d: y = 16'hfe00;
			16'hd88e: y = 16'hfe00;
			16'hd88f: y = 16'hfe00;
			16'hd890: y = 16'hfe00;
			16'hd891: y = 16'hfe00;
			16'hd892: y = 16'hfe00;
			16'hd893: y = 16'hfe00;
			16'hd894: y = 16'hfe00;
			16'hd895: y = 16'hfe00;
			16'hd896: y = 16'hfe00;
			16'hd897: y = 16'hfe00;
			16'hd898: y = 16'hfe00;
			16'hd899: y = 16'hfe00;
			16'hd89a: y = 16'hfe00;
			16'hd89b: y = 16'hfe00;
			16'hd89c: y = 16'hfe00;
			16'hd89d: y = 16'hfe00;
			16'hd89e: y = 16'hfe00;
			16'hd89f: y = 16'hfe00;
			16'hd8a0: y = 16'hfe00;
			16'hd8a1: y = 16'hfe00;
			16'hd8a2: y = 16'hfe00;
			16'hd8a3: y = 16'hfe00;
			16'hd8a4: y = 16'hfe00;
			16'hd8a5: y = 16'hfe00;
			16'hd8a6: y = 16'hfe00;
			16'hd8a7: y = 16'hfe00;
			16'hd8a8: y = 16'hfe00;
			16'hd8a9: y = 16'hfe00;
			16'hd8aa: y = 16'hfe00;
			16'hd8ab: y = 16'hfe00;
			16'hd8ac: y = 16'hfe00;
			16'hd8ad: y = 16'hfe00;
			16'hd8ae: y = 16'hfe00;
			16'hd8af: y = 16'hfe00;
			16'hd8b0: y = 16'hfe00;
			16'hd8b1: y = 16'hfe00;
			16'hd8b2: y = 16'hfe00;
			16'hd8b3: y = 16'hfe00;
			16'hd8b4: y = 16'hfe00;
			16'hd8b5: y = 16'hfe00;
			16'hd8b6: y = 16'hfe00;
			16'hd8b7: y = 16'hfe00;
			16'hd8b8: y = 16'hfe00;
			16'hd8b9: y = 16'hfe00;
			16'hd8ba: y = 16'hfe00;
			16'hd8bb: y = 16'hfe00;
			16'hd8bc: y = 16'hfe00;
			16'hd8bd: y = 16'hfe00;
			16'hd8be: y = 16'hfe00;
			16'hd8bf: y = 16'hfe00;
			16'hd8c0: y = 16'hfe00;
			16'hd8c1: y = 16'hfe00;
			16'hd8c2: y = 16'hfe00;
			16'hd8c3: y = 16'hfe00;
			16'hd8c4: y = 16'hfe00;
			16'hd8c5: y = 16'hfe00;
			16'hd8c6: y = 16'hfe00;
			16'hd8c7: y = 16'hfe00;
			16'hd8c8: y = 16'hfe00;
			16'hd8c9: y = 16'hfe00;
			16'hd8ca: y = 16'hfe00;
			16'hd8cb: y = 16'hfe00;
			16'hd8cc: y = 16'hfe00;
			16'hd8cd: y = 16'hfe00;
			16'hd8ce: y = 16'hfe00;
			16'hd8cf: y = 16'hfe00;
			16'hd8d0: y = 16'hfe00;
			16'hd8d1: y = 16'hfe00;
			16'hd8d2: y = 16'hfe00;
			16'hd8d3: y = 16'hfe00;
			16'hd8d4: y = 16'hfe00;
			16'hd8d5: y = 16'hfe00;
			16'hd8d6: y = 16'hfe00;
			16'hd8d7: y = 16'hfe00;
			16'hd8d8: y = 16'hfe00;
			16'hd8d9: y = 16'hfe00;
			16'hd8da: y = 16'hfe00;
			16'hd8db: y = 16'hfe00;
			16'hd8dc: y = 16'hfe00;
			16'hd8dd: y = 16'hfe00;
			16'hd8de: y = 16'hfe00;
			16'hd8df: y = 16'hfe00;
			16'hd8e0: y = 16'hfe00;
			16'hd8e1: y = 16'hfe00;
			16'hd8e2: y = 16'hfe00;
			16'hd8e3: y = 16'hfe00;
			16'hd8e4: y = 16'hfe00;
			16'hd8e5: y = 16'hfe00;
			16'hd8e6: y = 16'hfe00;
			16'hd8e7: y = 16'hfe00;
			16'hd8e8: y = 16'hfe00;
			16'hd8e9: y = 16'hfe00;
			16'hd8ea: y = 16'hfe00;
			16'hd8eb: y = 16'hfe00;
			16'hd8ec: y = 16'hfe00;
			16'hd8ed: y = 16'hfe00;
			16'hd8ee: y = 16'hfe00;
			16'hd8ef: y = 16'hfe00;
			16'hd8f0: y = 16'hfe00;
			16'hd8f1: y = 16'hfe00;
			16'hd8f2: y = 16'hfe00;
			16'hd8f3: y = 16'hfe00;
			16'hd8f4: y = 16'hfe00;
			16'hd8f5: y = 16'hfe00;
			16'hd8f6: y = 16'hfe00;
			16'hd8f7: y = 16'hfe00;
			16'hd8f8: y = 16'hfe00;
			16'hd8f9: y = 16'hfe00;
			16'hd8fa: y = 16'hfe00;
			16'hd8fb: y = 16'hfe00;
			16'hd8fc: y = 16'hfe00;
			16'hd8fd: y = 16'hfe00;
			16'hd8fe: y = 16'hfe00;
			16'hd8ff: y = 16'hfe00;
			16'hd900: y = 16'hfe00;
			16'hd901: y = 16'hfe00;
			16'hd902: y = 16'hfe00;
			16'hd903: y = 16'hfe00;
			16'hd904: y = 16'hfe00;
			16'hd905: y = 16'hfe00;
			16'hd906: y = 16'hfe00;
			16'hd907: y = 16'hfe00;
			16'hd908: y = 16'hfe00;
			16'hd909: y = 16'hfe00;
			16'hd90a: y = 16'hfe00;
			16'hd90b: y = 16'hfe00;
			16'hd90c: y = 16'hfe00;
			16'hd90d: y = 16'hfe00;
			16'hd90e: y = 16'hfe00;
			16'hd90f: y = 16'hfe00;
			16'hd910: y = 16'hfe00;
			16'hd911: y = 16'hfe00;
			16'hd912: y = 16'hfe00;
			16'hd913: y = 16'hfe00;
			16'hd914: y = 16'hfe00;
			16'hd915: y = 16'hfe00;
			16'hd916: y = 16'hfe00;
			16'hd917: y = 16'hfe00;
			16'hd918: y = 16'hfe00;
			16'hd919: y = 16'hfe00;
			16'hd91a: y = 16'hfe00;
			16'hd91b: y = 16'hfe00;
			16'hd91c: y = 16'hfe00;
			16'hd91d: y = 16'hfe00;
			16'hd91e: y = 16'hfe00;
			16'hd91f: y = 16'hfe00;
			16'hd920: y = 16'hfe00;
			16'hd921: y = 16'hfe00;
			16'hd922: y = 16'hfe00;
			16'hd923: y = 16'hfe00;
			16'hd924: y = 16'hfe00;
			16'hd925: y = 16'hfe00;
			16'hd926: y = 16'hfe00;
			16'hd927: y = 16'hfe00;
			16'hd928: y = 16'hfe00;
			16'hd929: y = 16'hfe00;
			16'hd92a: y = 16'hfe00;
			16'hd92b: y = 16'hfe00;
			16'hd92c: y = 16'hfe00;
			16'hd92d: y = 16'hfe00;
			16'hd92e: y = 16'hfe00;
			16'hd92f: y = 16'hfe00;
			16'hd930: y = 16'hfe00;
			16'hd931: y = 16'hfe00;
			16'hd932: y = 16'hfe00;
			16'hd933: y = 16'hfe00;
			16'hd934: y = 16'hfe00;
			16'hd935: y = 16'hfe00;
			16'hd936: y = 16'hfe00;
			16'hd937: y = 16'hfe00;
			16'hd938: y = 16'hfe00;
			16'hd939: y = 16'hfe00;
			16'hd93a: y = 16'hfe00;
			16'hd93b: y = 16'hfe00;
			16'hd93c: y = 16'hfe00;
			16'hd93d: y = 16'hfe00;
			16'hd93e: y = 16'hfe00;
			16'hd93f: y = 16'hfe00;
			16'hd940: y = 16'hfe00;
			16'hd941: y = 16'hfe00;
			16'hd942: y = 16'hfe00;
			16'hd943: y = 16'hfe00;
			16'hd944: y = 16'hfe00;
			16'hd945: y = 16'hfe00;
			16'hd946: y = 16'hfe00;
			16'hd947: y = 16'hfe00;
			16'hd948: y = 16'hfe00;
			16'hd949: y = 16'hfe00;
			16'hd94a: y = 16'hfe00;
			16'hd94b: y = 16'hfe00;
			16'hd94c: y = 16'hfe00;
			16'hd94d: y = 16'hfe00;
			16'hd94e: y = 16'hfe00;
			16'hd94f: y = 16'hfe00;
			16'hd950: y = 16'hfe00;
			16'hd951: y = 16'hfe00;
			16'hd952: y = 16'hfe00;
			16'hd953: y = 16'hfe00;
			16'hd954: y = 16'hfe00;
			16'hd955: y = 16'hfe00;
			16'hd956: y = 16'hfe00;
			16'hd957: y = 16'hfe00;
			16'hd958: y = 16'hfe00;
			16'hd959: y = 16'hfe00;
			16'hd95a: y = 16'hfe00;
			16'hd95b: y = 16'hfe00;
			16'hd95c: y = 16'hfe00;
			16'hd95d: y = 16'hfe00;
			16'hd95e: y = 16'hfe00;
			16'hd95f: y = 16'hfe00;
			16'hd960: y = 16'hfe00;
			16'hd961: y = 16'hfe00;
			16'hd962: y = 16'hfe00;
			16'hd963: y = 16'hfe00;
			16'hd964: y = 16'hfe00;
			16'hd965: y = 16'hfe00;
			16'hd966: y = 16'hfe00;
			16'hd967: y = 16'hfe00;
			16'hd968: y = 16'hfe00;
			16'hd969: y = 16'hfe00;
			16'hd96a: y = 16'hfe00;
			16'hd96b: y = 16'hfe00;
			16'hd96c: y = 16'hfe00;
			16'hd96d: y = 16'hfe00;
			16'hd96e: y = 16'hfe00;
			16'hd96f: y = 16'hfe00;
			16'hd970: y = 16'hfe00;
			16'hd971: y = 16'hfe00;
			16'hd972: y = 16'hfe00;
			16'hd973: y = 16'hfe00;
			16'hd974: y = 16'hfe00;
			16'hd975: y = 16'hfe00;
			16'hd976: y = 16'hfe00;
			16'hd977: y = 16'hfe00;
			16'hd978: y = 16'hfe00;
			16'hd979: y = 16'hfe00;
			16'hd97a: y = 16'hfe00;
			16'hd97b: y = 16'hfe00;
			16'hd97c: y = 16'hfe00;
			16'hd97d: y = 16'hfe00;
			16'hd97e: y = 16'hfe00;
			16'hd97f: y = 16'hfe00;
			16'hd980: y = 16'hfe00;
			16'hd981: y = 16'hfe00;
			16'hd982: y = 16'hfe00;
			16'hd983: y = 16'hfe00;
			16'hd984: y = 16'hfe00;
			16'hd985: y = 16'hfe00;
			16'hd986: y = 16'hfe00;
			16'hd987: y = 16'hfe00;
			16'hd988: y = 16'hfe00;
			16'hd989: y = 16'hfe00;
			16'hd98a: y = 16'hfe00;
			16'hd98b: y = 16'hfe00;
			16'hd98c: y = 16'hfe00;
			16'hd98d: y = 16'hfe00;
			16'hd98e: y = 16'hfe00;
			16'hd98f: y = 16'hfe00;
			16'hd990: y = 16'hfe00;
			16'hd991: y = 16'hfe00;
			16'hd992: y = 16'hfe00;
			16'hd993: y = 16'hfe00;
			16'hd994: y = 16'hfe00;
			16'hd995: y = 16'hfe00;
			16'hd996: y = 16'hfe00;
			16'hd997: y = 16'hfe00;
			16'hd998: y = 16'hfe00;
			16'hd999: y = 16'hfe00;
			16'hd99a: y = 16'hfe00;
			16'hd99b: y = 16'hfe00;
			16'hd99c: y = 16'hfe00;
			16'hd99d: y = 16'hfe00;
			16'hd99e: y = 16'hfe00;
			16'hd99f: y = 16'hfe00;
			16'hd9a0: y = 16'hfe00;
			16'hd9a1: y = 16'hfe00;
			16'hd9a2: y = 16'hfe00;
			16'hd9a3: y = 16'hfe00;
			16'hd9a4: y = 16'hfe00;
			16'hd9a5: y = 16'hfe00;
			16'hd9a6: y = 16'hfe00;
			16'hd9a7: y = 16'hfe00;
			16'hd9a8: y = 16'hfe00;
			16'hd9a9: y = 16'hfe00;
			16'hd9aa: y = 16'hfe00;
			16'hd9ab: y = 16'hfe00;
			16'hd9ac: y = 16'hfe00;
			16'hd9ad: y = 16'hfe00;
			16'hd9ae: y = 16'hfe00;
			16'hd9af: y = 16'hfe00;
			16'hd9b0: y = 16'hfe00;
			16'hd9b1: y = 16'hfe00;
			16'hd9b2: y = 16'hfe00;
			16'hd9b3: y = 16'hfe00;
			16'hd9b4: y = 16'hfe00;
			16'hd9b5: y = 16'hfe00;
			16'hd9b6: y = 16'hfe00;
			16'hd9b7: y = 16'hfe00;
			16'hd9b8: y = 16'hfe00;
			16'hd9b9: y = 16'hfe00;
			16'hd9ba: y = 16'hfe00;
			16'hd9bb: y = 16'hfe00;
			16'hd9bc: y = 16'hfe00;
			16'hd9bd: y = 16'hfe00;
			16'hd9be: y = 16'hfe00;
			16'hd9bf: y = 16'hfe00;
			16'hd9c0: y = 16'hfe00;
			16'hd9c1: y = 16'hfe00;
			16'hd9c2: y = 16'hfe00;
			16'hd9c3: y = 16'hfe00;
			16'hd9c4: y = 16'hfe00;
			16'hd9c5: y = 16'hfe00;
			16'hd9c6: y = 16'hfe00;
			16'hd9c7: y = 16'hfe00;
			16'hd9c8: y = 16'hfe00;
			16'hd9c9: y = 16'hfe00;
			16'hd9ca: y = 16'hfe00;
			16'hd9cb: y = 16'hfe00;
			16'hd9cc: y = 16'hfe00;
			16'hd9cd: y = 16'hfe00;
			16'hd9ce: y = 16'hfe00;
			16'hd9cf: y = 16'hfe00;
			16'hd9d0: y = 16'hfe00;
			16'hd9d1: y = 16'hfe00;
			16'hd9d2: y = 16'hfe00;
			16'hd9d3: y = 16'hfe00;
			16'hd9d4: y = 16'hfe00;
			16'hd9d5: y = 16'hfe00;
			16'hd9d6: y = 16'hfe00;
			16'hd9d7: y = 16'hfe00;
			16'hd9d8: y = 16'hfe00;
			16'hd9d9: y = 16'hfe00;
			16'hd9da: y = 16'hfe00;
			16'hd9db: y = 16'hfe00;
			16'hd9dc: y = 16'hfe00;
			16'hd9dd: y = 16'hfe00;
			16'hd9de: y = 16'hfe00;
			16'hd9df: y = 16'hfe00;
			16'hd9e0: y = 16'hfe00;
			16'hd9e1: y = 16'hfe00;
			16'hd9e2: y = 16'hfe00;
			16'hd9e3: y = 16'hfe00;
			16'hd9e4: y = 16'hfe00;
			16'hd9e5: y = 16'hfe00;
			16'hd9e6: y = 16'hfe00;
			16'hd9e7: y = 16'hfe00;
			16'hd9e8: y = 16'hfe00;
			16'hd9e9: y = 16'hfe00;
			16'hd9ea: y = 16'hfe00;
			16'hd9eb: y = 16'hfe00;
			16'hd9ec: y = 16'hfe00;
			16'hd9ed: y = 16'hfe00;
			16'hd9ee: y = 16'hfe00;
			16'hd9ef: y = 16'hfe00;
			16'hd9f0: y = 16'hfe00;
			16'hd9f1: y = 16'hfe00;
			16'hd9f2: y = 16'hfe00;
			16'hd9f3: y = 16'hfe00;
			16'hd9f4: y = 16'hfe00;
			16'hd9f5: y = 16'hfe00;
			16'hd9f6: y = 16'hfe00;
			16'hd9f7: y = 16'hfe00;
			16'hd9f8: y = 16'hfe00;
			16'hd9f9: y = 16'hfe00;
			16'hd9fa: y = 16'hfe00;
			16'hd9fb: y = 16'hfe00;
			16'hd9fc: y = 16'hfe00;
			16'hd9fd: y = 16'hfe00;
			16'hd9fe: y = 16'hfe00;
			16'hd9ff: y = 16'hfe00;
			16'hda00: y = 16'hfe00;
			16'hda01: y = 16'hfe00;
			16'hda02: y = 16'hfe00;
			16'hda03: y = 16'hfe00;
			16'hda04: y = 16'hfe00;
			16'hda05: y = 16'hfe00;
			16'hda06: y = 16'hfe00;
			16'hda07: y = 16'hfe00;
			16'hda08: y = 16'hfe00;
			16'hda09: y = 16'hfe00;
			16'hda0a: y = 16'hfe00;
			16'hda0b: y = 16'hfe00;
			16'hda0c: y = 16'hfe00;
			16'hda0d: y = 16'hfe00;
			16'hda0e: y = 16'hfe00;
			16'hda0f: y = 16'hfe00;
			16'hda10: y = 16'hfe00;
			16'hda11: y = 16'hfe00;
			16'hda12: y = 16'hfe00;
			16'hda13: y = 16'hfe00;
			16'hda14: y = 16'hfe00;
			16'hda15: y = 16'hfe00;
			16'hda16: y = 16'hfe00;
			16'hda17: y = 16'hfe00;
			16'hda18: y = 16'hfe00;
			16'hda19: y = 16'hfe00;
			16'hda1a: y = 16'hfe00;
			16'hda1b: y = 16'hfe00;
			16'hda1c: y = 16'hfe00;
			16'hda1d: y = 16'hfe00;
			16'hda1e: y = 16'hfe00;
			16'hda1f: y = 16'hfe00;
			16'hda20: y = 16'hfe00;
			16'hda21: y = 16'hfe00;
			16'hda22: y = 16'hfe00;
			16'hda23: y = 16'hfe00;
			16'hda24: y = 16'hfe00;
			16'hda25: y = 16'hfe00;
			16'hda26: y = 16'hfe00;
			16'hda27: y = 16'hfe00;
			16'hda28: y = 16'hfe00;
			16'hda29: y = 16'hfe00;
			16'hda2a: y = 16'hfe00;
			16'hda2b: y = 16'hfe00;
			16'hda2c: y = 16'hfe00;
			16'hda2d: y = 16'hfe00;
			16'hda2e: y = 16'hfe00;
			16'hda2f: y = 16'hfe00;
			16'hda30: y = 16'hfe00;
			16'hda31: y = 16'hfe00;
			16'hda32: y = 16'hfe00;
			16'hda33: y = 16'hfe00;
			16'hda34: y = 16'hfe00;
			16'hda35: y = 16'hfe00;
			16'hda36: y = 16'hfe00;
			16'hda37: y = 16'hfe00;
			16'hda38: y = 16'hfe00;
			16'hda39: y = 16'hfe00;
			16'hda3a: y = 16'hfe00;
			16'hda3b: y = 16'hfe00;
			16'hda3c: y = 16'hfe00;
			16'hda3d: y = 16'hfe00;
			16'hda3e: y = 16'hfe00;
			16'hda3f: y = 16'hfe00;
			16'hda40: y = 16'hfe00;
			16'hda41: y = 16'hfe00;
			16'hda42: y = 16'hfe00;
			16'hda43: y = 16'hfe00;
			16'hda44: y = 16'hfe00;
			16'hda45: y = 16'hfe00;
			16'hda46: y = 16'hfe00;
			16'hda47: y = 16'hfe00;
			16'hda48: y = 16'hfe00;
			16'hda49: y = 16'hfe00;
			16'hda4a: y = 16'hfe00;
			16'hda4b: y = 16'hfe00;
			16'hda4c: y = 16'hfe00;
			16'hda4d: y = 16'hfe00;
			16'hda4e: y = 16'hfe00;
			16'hda4f: y = 16'hfe00;
			16'hda50: y = 16'hfe00;
			16'hda51: y = 16'hfe00;
			16'hda52: y = 16'hfe00;
			16'hda53: y = 16'hfe00;
			16'hda54: y = 16'hfe00;
			16'hda55: y = 16'hfe00;
			16'hda56: y = 16'hfe00;
			16'hda57: y = 16'hfe00;
			16'hda58: y = 16'hfe00;
			16'hda59: y = 16'hfe00;
			16'hda5a: y = 16'hfe00;
			16'hda5b: y = 16'hfe00;
			16'hda5c: y = 16'hfe00;
			16'hda5d: y = 16'hfe00;
			16'hda5e: y = 16'hfe00;
			16'hda5f: y = 16'hfe00;
			16'hda60: y = 16'hfe00;
			16'hda61: y = 16'hfe00;
			16'hda62: y = 16'hfe00;
			16'hda63: y = 16'hfe00;
			16'hda64: y = 16'hfe00;
			16'hda65: y = 16'hfe00;
			16'hda66: y = 16'hfe00;
			16'hda67: y = 16'hfe00;
			16'hda68: y = 16'hfe00;
			16'hda69: y = 16'hfe00;
			16'hda6a: y = 16'hfe00;
			16'hda6b: y = 16'hfe00;
			16'hda6c: y = 16'hfe00;
			16'hda6d: y = 16'hfe00;
			16'hda6e: y = 16'hfe00;
			16'hda6f: y = 16'hfe00;
			16'hda70: y = 16'hfe00;
			16'hda71: y = 16'hfe00;
			16'hda72: y = 16'hfe00;
			16'hda73: y = 16'hfe00;
			16'hda74: y = 16'hfe00;
			16'hda75: y = 16'hfe00;
			16'hda76: y = 16'hfe00;
			16'hda77: y = 16'hfe00;
			16'hda78: y = 16'hfe00;
			16'hda79: y = 16'hfe00;
			16'hda7a: y = 16'hfe00;
			16'hda7b: y = 16'hfe00;
			16'hda7c: y = 16'hfe00;
			16'hda7d: y = 16'hfe00;
			16'hda7e: y = 16'hfe00;
			16'hda7f: y = 16'hfe00;
			16'hda80: y = 16'hfe00;
			16'hda81: y = 16'hfe00;
			16'hda82: y = 16'hfe00;
			16'hda83: y = 16'hfe00;
			16'hda84: y = 16'hfe00;
			16'hda85: y = 16'hfe00;
			16'hda86: y = 16'hfe00;
			16'hda87: y = 16'hfe00;
			16'hda88: y = 16'hfe00;
			16'hda89: y = 16'hfe00;
			16'hda8a: y = 16'hfe00;
			16'hda8b: y = 16'hfe00;
			16'hda8c: y = 16'hfe00;
			16'hda8d: y = 16'hfe00;
			16'hda8e: y = 16'hfe00;
			16'hda8f: y = 16'hfe00;
			16'hda90: y = 16'hfe00;
			16'hda91: y = 16'hfe00;
			16'hda92: y = 16'hfe01;
			16'hda93: y = 16'hfe01;
			16'hda94: y = 16'hfe01;
			16'hda95: y = 16'hfe01;
			16'hda96: y = 16'hfe01;
			16'hda97: y = 16'hfe01;
			16'hda98: y = 16'hfe01;
			16'hda99: y = 16'hfe01;
			16'hda9a: y = 16'hfe01;
			16'hda9b: y = 16'hfe01;
			16'hda9c: y = 16'hfe01;
			16'hda9d: y = 16'hfe01;
			16'hda9e: y = 16'hfe01;
			16'hda9f: y = 16'hfe01;
			16'hdaa0: y = 16'hfe01;
			16'hdaa1: y = 16'hfe01;
			16'hdaa2: y = 16'hfe01;
			16'hdaa3: y = 16'hfe01;
			16'hdaa4: y = 16'hfe01;
			16'hdaa5: y = 16'hfe01;
			16'hdaa6: y = 16'hfe01;
			16'hdaa7: y = 16'hfe01;
			16'hdaa8: y = 16'hfe01;
			16'hdaa9: y = 16'hfe01;
			16'hdaaa: y = 16'hfe01;
			16'hdaab: y = 16'hfe01;
			16'hdaac: y = 16'hfe01;
			16'hdaad: y = 16'hfe01;
			16'hdaae: y = 16'hfe01;
			16'hdaaf: y = 16'hfe01;
			16'hdab0: y = 16'hfe01;
			16'hdab1: y = 16'hfe01;
			16'hdab2: y = 16'hfe01;
			16'hdab3: y = 16'hfe01;
			16'hdab4: y = 16'hfe01;
			16'hdab5: y = 16'hfe01;
			16'hdab6: y = 16'hfe01;
			16'hdab7: y = 16'hfe01;
			16'hdab8: y = 16'hfe01;
			16'hdab9: y = 16'hfe01;
			16'hdaba: y = 16'hfe01;
			16'hdabb: y = 16'hfe01;
			16'hdabc: y = 16'hfe01;
			16'hdabd: y = 16'hfe01;
			16'hdabe: y = 16'hfe01;
			16'hdabf: y = 16'hfe01;
			16'hdac0: y = 16'hfe01;
			16'hdac1: y = 16'hfe01;
			16'hdac2: y = 16'hfe01;
			16'hdac3: y = 16'hfe01;
			16'hdac4: y = 16'hfe01;
			16'hdac5: y = 16'hfe01;
			16'hdac6: y = 16'hfe01;
			16'hdac7: y = 16'hfe01;
			16'hdac8: y = 16'hfe01;
			16'hdac9: y = 16'hfe01;
			16'hdaca: y = 16'hfe01;
			16'hdacb: y = 16'hfe01;
			16'hdacc: y = 16'hfe01;
			16'hdacd: y = 16'hfe01;
			16'hdace: y = 16'hfe01;
			16'hdacf: y = 16'hfe01;
			16'hdad0: y = 16'hfe01;
			16'hdad1: y = 16'hfe01;
			16'hdad2: y = 16'hfe01;
			16'hdad3: y = 16'hfe01;
			16'hdad4: y = 16'hfe01;
			16'hdad5: y = 16'hfe01;
			16'hdad6: y = 16'hfe01;
			16'hdad7: y = 16'hfe01;
			16'hdad8: y = 16'hfe01;
			16'hdad9: y = 16'hfe01;
			16'hdada: y = 16'hfe01;
			16'hdadb: y = 16'hfe01;
			16'hdadc: y = 16'hfe01;
			16'hdadd: y = 16'hfe01;
			16'hdade: y = 16'hfe01;
			16'hdadf: y = 16'hfe01;
			16'hdae0: y = 16'hfe01;
			16'hdae1: y = 16'hfe01;
			16'hdae2: y = 16'hfe01;
			16'hdae3: y = 16'hfe01;
			16'hdae4: y = 16'hfe01;
			16'hdae5: y = 16'hfe01;
			16'hdae6: y = 16'hfe01;
			16'hdae7: y = 16'hfe01;
			16'hdae8: y = 16'hfe01;
			16'hdae9: y = 16'hfe01;
			16'hdaea: y = 16'hfe01;
			16'hdaeb: y = 16'hfe01;
			16'hdaec: y = 16'hfe01;
			16'hdaed: y = 16'hfe01;
			16'hdaee: y = 16'hfe01;
			16'hdaef: y = 16'hfe01;
			16'hdaf0: y = 16'hfe01;
			16'hdaf1: y = 16'hfe01;
			16'hdaf2: y = 16'hfe01;
			16'hdaf3: y = 16'hfe01;
			16'hdaf4: y = 16'hfe01;
			16'hdaf5: y = 16'hfe01;
			16'hdaf6: y = 16'hfe01;
			16'hdaf7: y = 16'hfe01;
			16'hdaf8: y = 16'hfe01;
			16'hdaf9: y = 16'hfe01;
			16'hdafa: y = 16'hfe01;
			16'hdafb: y = 16'hfe01;
			16'hdafc: y = 16'hfe01;
			16'hdafd: y = 16'hfe01;
			16'hdafe: y = 16'hfe01;
			16'hdaff: y = 16'hfe01;
			16'hdb00: y = 16'hfe01;
			16'hdb01: y = 16'hfe01;
			16'hdb02: y = 16'hfe01;
			16'hdb03: y = 16'hfe01;
			16'hdb04: y = 16'hfe01;
			16'hdb05: y = 16'hfe01;
			16'hdb06: y = 16'hfe01;
			16'hdb07: y = 16'hfe01;
			16'hdb08: y = 16'hfe01;
			16'hdb09: y = 16'hfe01;
			16'hdb0a: y = 16'hfe01;
			16'hdb0b: y = 16'hfe01;
			16'hdb0c: y = 16'hfe01;
			16'hdb0d: y = 16'hfe01;
			16'hdb0e: y = 16'hfe01;
			16'hdb0f: y = 16'hfe01;
			16'hdb10: y = 16'hfe01;
			16'hdb11: y = 16'hfe01;
			16'hdb12: y = 16'hfe01;
			16'hdb13: y = 16'hfe01;
			16'hdb14: y = 16'hfe01;
			16'hdb15: y = 16'hfe01;
			16'hdb16: y = 16'hfe01;
			16'hdb17: y = 16'hfe01;
			16'hdb18: y = 16'hfe01;
			16'hdb19: y = 16'hfe01;
			16'hdb1a: y = 16'hfe01;
			16'hdb1b: y = 16'hfe01;
			16'hdb1c: y = 16'hfe01;
			16'hdb1d: y = 16'hfe01;
			16'hdb1e: y = 16'hfe01;
			16'hdb1f: y = 16'hfe01;
			16'hdb20: y = 16'hfe01;
			16'hdb21: y = 16'hfe01;
			16'hdb22: y = 16'hfe01;
			16'hdb23: y = 16'hfe01;
			16'hdb24: y = 16'hfe01;
			16'hdb25: y = 16'hfe01;
			16'hdb26: y = 16'hfe01;
			16'hdb27: y = 16'hfe01;
			16'hdb28: y = 16'hfe01;
			16'hdb29: y = 16'hfe01;
			16'hdb2a: y = 16'hfe01;
			16'hdb2b: y = 16'hfe01;
			16'hdb2c: y = 16'hfe01;
			16'hdb2d: y = 16'hfe01;
			16'hdb2e: y = 16'hfe01;
			16'hdb2f: y = 16'hfe01;
			16'hdb30: y = 16'hfe01;
			16'hdb31: y = 16'hfe01;
			16'hdb32: y = 16'hfe01;
			16'hdb33: y = 16'hfe01;
			16'hdb34: y = 16'hfe01;
			16'hdb35: y = 16'hfe01;
			16'hdb36: y = 16'hfe01;
			16'hdb37: y = 16'hfe01;
			16'hdb38: y = 16'hfe01;
			16'hdb39: y = 16'hfe01;
			16'hdb3a: y = 16'hfe01;
			16'hdb3b: y = 16'hfe01;
			16'hdb3c: y = 16'hfe01;
			16'hdb3d: y = 16'hfe01;
			16'hdb3e: y = 16'hfe01;
			16'hdb3f: y = 16'hfe01;
			16'hdb40: y = 16'hfe01;
			16'hdb41: y = 16'hfe01;
			16'hdb42: y = 16'hfe01;
			16'hdb43: y = 16'hfe01;
			16'hdb44: y = 16'hfe01;
			16'hdb45: y = 16'hfe01;
			16'hdb46: y = 16'hfe01;
			16'hdb47: y = 16'hfe01;
			16'hdb48: y = 16'hfe01;
			16'hdb49: y = 16'hfe01;
			16'hdb4a: y = 16'hfe01;
			16'hdb4b: y = 16'hfe01;
			16'hdb4c: y = 16'hfe01;
			16'hdb4d: y = 16'hfe01;
			16'hdb4e: y = 16'hfe01;
			16'hdb4f: y = 16'hfe01;
			16'hdb50: y = 16'hfe01;
			16'hdb51: y = 16'hfe01;
			16'hdb52: y = 16'hfe01;
			16'hdb53: y = 16'hfe01;
			16'hdb54: y = 16'hfe01;
			16'hdb55: y = 16'hfe01;
			16'hdb56: y = 16'hfe01;
			16'hdb57: y = 16'hfe01;
			16'hdb58: y = 16'hfe01;
			16'hdb59: y = 16'hfe01;
			16'hdb5a: y = 16'hfe01;
			16'hdb5b: y = 16'hfe01;
			16'hdb5c: y = 16'hfe01;
			16'hdb5d: y = 16'hfe01;
			16'hdb5e: y = 16'hfe01;
			16'hdb5f: y = 16'hfe01;
			16'hdb60: y = 16'hfe01;
			16'hdb61: y = 16'hfe01;
			16'hdb62: y = 16'hfe01;
			16'hdb63: y = 16'hfe01;
			16'hdb64: y = 16'hfe01;
			16'hdb65: y = 16'hfe01;
			16'hdb66: y = 16'hfe01;
			16'hdb67: y = 16'hfe01;
			16'hdb68: y = 16'hfe01;
			16'hdb69: y = 16'hfe01;
			16'hdb6a: y = 16'hfe01;
			16'hdb6b: y = 16'hfe01;
			16'hdb6c: y = 16'hfe01;
			16'hdb6d: y = 16'hfe01;
			16'hdb6e: y = 16'hfe01;
			16'hdb6f: y = 16'hfe01;
			16'hdb70: y = 16'hfe01;
			16'hdb71: y = 16'hfe01;
			16'hdb72: y = 16'hfe01;
			16'hdb73: y = 16'hfe01;
			16'hdb74: y = 16'hfe01;
			16'hdb75: y = 16'hfe01;
			16'hdb76: y = 16'hfe01;
			16'hdb77: y = 16'hfe01;
			16'hdb78: y = 16'hfe01;
			16'hdb79: y = 16'hfe01;
			16'hdb7a: y = 16'hfe01;
			16'hdb7b: y = 16'hfe01;
			16'hdb7c: y = 16'hfe01;
			16'hdb7d: y = 16'hfe01;
			16'hdb7e: y = 16'hfe01;
			16'hdb7f: y = 16'hfe01;
			16'hdb80: y = 16'hfe01;
			16'hdb81: y = 16'hfe01;
			16'hdb82: y = 16'hfe01;
			16'hdb83: y = 16'hfe01;
			16'hdb84: y = 16'hfe01;
			16'hdb85: y = 16'hfe01;
			16'hdb86: y = 16'hfe01;
			16'hdb87: y = 16'hfe01;
			16'hdb88: y = 16'hfe01;
			16'hdb89: y = 16'hfe01;
			16'hdb8a: y = 16'hfe01;
			16'hdb8b: y = 16'hfe01;
			16'hdb8c: y = 16'hfe01;
			16'hdb8d: y = 16'hfe01;
			16'hdb8e: y = 16'hfe01;
			16'hdb8f: y = 16'hfe01;
			16'hdb90: y = 16'hfe01;
			16'hdb91: y = 16'hfe01;
			16'hdb92: y = 16'hfe01;
			16'hdb93: y = 16'hfe01;
			16'hdb94: y = 16'hfe01;
			16'hdb95: y = 16'hfe01;
			16'hdb96: y = 16'hfe01;
			16'hdb97: y = 16'hfe01;
			16'hdb98: y = 16'hfe01;
			16'hdb99: y = 16'hfe01;
			16'hdb9a: y = 16'hfe01;
			16'hdb9b: y = 16'hfe01;
			16'hdb9c: y = 16'hfe01;
			16'hdb9d: y = 16'hfe01;
			16'hdb9e: y = 16'hfe01;
			16'hdb9f: y = 16'hfe01;
			16'hdba0: y = 16'hfe01;
			16'hdba1: y = 16'hfe01;
			16'hdba2: y = 16'hfe01;
			16'hdba3: y = 16'hfe01;
			16'hdba4: y = 16'hfe01;
			16'hdba5: y = 16'hfe01;
			16'hdba6: y = 16'hfe01;
			16'hdba7: y = 16'hfe01;
			16'hdba8: y = 16'hfe01;
			16'hdba9: y = 16'hfe01;
			16'hdbaa: y = 16'hfe01;
			16'hdbab: y = 16'hfe01;
			16'hdbac: y = 16'hfe01;
			16'hdbad: y = 16'hfe01;
			16'hdbae: y = 16'hfe01;
			16'hdbaf: y = 16'hfe01;
			16'hdbb0: y = 16'hfe01;
			16'hdbb1: y = 16'hfe01;
			16'hdbb2: y = 16'hfe01;
			16'hdbb3: y = 16'hfe01;
			16'hdbb4: y = 16'hfe01;
			16'hdbb5: y = 16'hfe01;
			16'hdbb6: y = 16'hfe01;
			16'hdbb7: y = 16'hfe01;
			16'hdbb8: y = 16'hfe01;
			16'hdbb9: y = 16'hfe01;
			16'hdbba: y = 16'hfe01;
			16'hdbbb: y = 16'hfe01;
			16'hdbbc: y = 16'hfe01;
			16'hdbbd: y = 16'hfe01;
			16'hdbbe: y = 16'hfe01;
			16'hdbbf: y = 16'hfe01;
			16'hdbc0: y = 16'hfe01;
			16'hdbc1: y = 16'hfe01;
			16'hdbc2: y = 16'hfe01;
			16'hdbc3: y = 16'hfe01;
			16'hdbc4: y = 16'hfe01;
			16'hdbc5: y = 16'hfe01;
			16'hdbc6: y = 16'hfe01;
			16'hdbc7: y = 16'hfe01;
			16'hdbc8: y = 16'hfe01;
			16'hdbc9: y = 16'hfe01;
			16'hdbca: y = 16'hfe01;
			16'hdbcb: y = 16'hfe01;
			16'hdbcc: y = 16'hfe01;
			16'hdbcd: y = 16'hfe01;
			16'hdbce: y = 16'hfe01;
			16'hdbcf: y = 16'hfe01;
			16'hdbd0: y = 16'hfe01;
			16'hdbd1: y = 16'hfe01;
			16'hdbd2: y = 16'hfe01;
			16'hdbd3: y = 16'hfe01;
			16'hdbd4: y = 16'hfe01;
			16'hdbd5: y = 16'hfe01;
			16'hdbd6: y = 16'hfe01;
			16'hdbd7: y = 16'hfe01;
			16'hdbd8: y = 16'hfe01;
			16'hdbd9: y = 16'hfe01;
			16'hdbda: y = 16'hfe01;
			16'hdbdb: y = 16'hfe01;
			16'hdbdc: y = 16'hfe01;
			16'hdbdd: y = 16'hfe01;
			16'hdbde: y = 16'hfe01;
			16'hdbdf: y = 16'hfe01;
			16'hdbe0: y = 16'hfe01;
			16'hdbe1: y = 16'hfe01;
			16'hdbe2: y = 16'hfe01;
			16'hdbe3: y = 16'hfe01;
			16'hdbe4: y = 16'hfe01;
			16'hdbe5: y = 16'hfe01;
			16'hdbe6: y = 16'hfe01;
			16'hdbe7: y = 16'hfe01;
			16'hdbe8: y = 16'hfe01;
			16'hdbe9: y = 16'hfe01;
			16'hdbea: y = 16'hfe01;
			16'hdbeb: y = 16'hfe01;
			16'hdbec: y = 16'hfe01;
			16'hdbed: y = 16'hfe01;
			16'hdbee: y = 16'hfe01;
			16'hdbef: y = 16'hfe01;
			16'hdbf0: y = 16'hfe01;
			16'hdbf1: y = 16'hfe01;
			16'hdbf2: y = 16'hfe01;
			16'hdbf3: y = 16'hfe01;
			16'hdbf4: y = 16'hfe01;
			16'hdbf5: y = 16'hfe01;
			16'hdbf6: y = 16'hfe01;
			16'hdbf7: y = 16'hfe01;
			16'hdbf8: y = 16'hfe01;
			16'hdbf9: y = 16'hfe01;
			16'hdbfa: y = 16'hfe01;
			16'hdbfb: y = 16'hfe01;
			16'hdbfc: y = 16'hfe01;
			16'hdbfd: y = 16'hfe01;
			16'hdbfe: y = 16'hfe01;
			16'hdbff: y = 16'hfe01;
			16'hdc00: y = 16'hfe01;
			16'hdc01: y = 16'hfe01;
			16'hdc02: y = 16'hfe01;
			16'hdc03: y = 16'hfe01;
			16'hdc04: y = 16'hfe01;
			16'hdc05: y = 16'hfe01;
			16'hdc06: y = 16'hfe01;
			16'hdc07: y = 16'hfe01;
			16'hdc08: y = 16'hfe01;
			16'hdc09: y = 16'hfe01;
			16'hdc0a: y = 16'hfe01;
			16'hdc0b: y = 16'hfe01;
			16'hdc0c: y = 16'hfe01;
			16'hdc0d: y = 16'hfe01;
			16'hdc0e: y = 16'hfe01;
			16'hdc0f: y = 16'hfe01;
			16'hdc10: y = 16'hfe01;
			16'hdc11: y = 16'hfe01;
			16'hdc12: y = 16'hfe01;
			16'hdc13: y = 16'hfe01;
			16'hdc14: y = 16'hfe01;
			16'hdc15: y = 16'hfe01;
			16'hdc16: y = 16'hfe01;
			16'hdc17: y = 16'hfe01;
			16'hdc18: y = 16'hfe01;
			16'hdc19: y = 16'hfe01;
			16'hdc1a: y = 16'hfe01;
			16'hdc1b: y = 16'hfe01;
			16'hdc1c: y = 16'hfe01;
			16'hdc1d: y = 16'hfe01;
			16'hdc1e: y = 16'hfe01;
			16'hdc1f: y = 16'hfe01;
			16'hdc20: y = 16'hfe01;
			16'hdc21: y = 16'hfe01;
			16'hdc22: y = 16'hfe01;
			16'hdc23: y = 16'hfe01;
			16'hdc24: y = 16'hfe01;
			16'hdc25: y = 16'hfe01;
			16'hdc26: y = 16'hfe01;
			16'hdc27: y = 16'hfe01;
			16'hdc28: y = 16'hfe01;
			16'hdc29: y = 16'hfe01;
			16'hdc2a: y = 16'hfe01;
			16'hdc2b: y = 16'hfe01;
			16'hdc2c: y = 16'hfe01;
			16'hdc2d: y = 16'hfe01;
			16'hdc2e: y = 16'hfe01;
			16'hdc2f: y = 16'hfe01;
			16'hdc30: y = 16'hfe01;
			16'hdc31: y = 16'hfe01;
			16'hdc32: y = 16'hfe01;
			16'hdc33: y = 16'hfe01;
			16'hdc34: y = 16'hfe01;
			16'hdc35: y = 16'hfe01;
			16'hdc36: y = 16'hfe01;
			16'hdc37: y = 16'hfe01;
			16'hdc38: y = 16'hfe01;
			16'hdc39: y = 16'hfe01;
			16'hdc3a: y = 16'hfe01;
			16'hdc3b: y = 16'hfe01;
			16'hdc3c: y = 16'hfe01;
			16'hdc3d: y = 16'hfe01;
			16'hdc3e: y = 16'hfe01;
			16'hdc3f: y = 16'hfe01;
			16'hdc40: y = 16'hfe01;
			16'hdc41: y = 16'hfe01;
			16'hdc42: y = 16'hfe01;
			16'hdc43: y = 16'hfe01;
			16'hdc44: y = 16'hfe01;
			16'hdc45: y = 16'hfe01;
			16'hdc46: y = 16'hfe01;
			16'hdc47: y = 16'hfe01;
			16'hdc48: y = 16'hfe01;
			16'hdc49: y = 16'hfe01;
			16'hdc4a: y = 16'hfe01;
			16'hdc4b: y = 16'hfe01;
			16'hdc4c: y = 16'hfe01;
			16'hdc4d: y = 16'hfe01;
			16'hdc4e: y = 16'hfe01;
			16'hdc4f: y = 16'hfe01;
			16'hdc50: y = 16'hfe01;
			16'hdc51: y = 16'hfe01;
			16'hdc52: y = 16'hfe01;
			16'hdc53: y = 16'hfe01;
			16'hdc54: y = 16'hfe01;
			16'hdc55: y = 16'hfe01;
			16'hdc56: y = 16'hfe01;
			16'hdc57: y = 16'hfe01;
			16'hdc58: y = 16'hfe01;
			16'hdc59: y = 16'hfe01;
			16'hdc5a: y = 16'hfe01;
			16'hdc5b: y = 16'hfe01;
			16'hdc5c: y = 16'hfe01;
			16'hdc5d: y = 16'hfe01;
			16'hdc5e: y = 16'hfe01;
			16'hdc5f: y = 16'hfe01;
			16'hdc60: y = 16'hfe01;
			16'hdc61: y = 16'hfe01;
			16'hdc62: y = 16'hfe01;
			16'hdc63: y = 16'hfe01;
			16'hdc64: y = 16'hfe01;
			16'hdc65: y = 16'hfe01;
			16'hdc66: y = 16'hfe01;
			16'hdc67: y = 16'hfe01;
			16'hdc68: y = 16'hfe01;
			16'hdc69: y = 16'hfe01;
			16'hdc6a: y = 16'hfe01;
			16'hdc6b: y = 16'hfe01;
			16'hdc6c: y = 16'hfe01;
			16'hdc6d: y = 16'hfe01;
			16'hdc6e: y = 16'hfe01;
			16'hdc6f: y = 16'hfe01;
			16'hdc70: y = 16'hfe01;
			16'hdc71: y = 16'hfe01;
			16'hdc72: y = 16'hfe01;
			16'hdc73: y = 16'hfe01;
			16'hdc74: y = 16'hfe01;
			16'hdc75: y = 16'hfe01;
			16'hdc76: y = 16'hfe01;
			16'hdc77: y = 16'hfe01;
			16'hdc78: y = 16'hfe01;
			16'hdc79: y = 16'hfe01;
			16'hdc7a: y = 16'hfe01;
			16'hdc7b: y = 16'hfe01;
			16'hdc7c: y = 16'hfe01;
			16'hdc7d: y = 16'hfe01;
			16'hdc7e: y = 16'hfe01;
			16'hdc7f: y = 16'hfe01;
			16'hdc80: y = 16'hfe01;
			16'hdc81: y = 16'hfe01;
			16'hdc82: y = 16'hfe01;
			16'hdc83: y = 16'hfe01;
			16'hdc84: y = 16'hfe01;
			16'hdc85: y = 16'hfe01;
			16'hdc86: y = 16'hfe01;
			16'hdc87: y = 16'hfe01;
			16'hdc88: y = 16'hfe01;
			16'hdc89: y = 16'hfe01;
			16'hdc8a: y = 16'hfe01;
			16'hdc8b: y = 16'hfe01;
			16'hdc8c: y = 16'hfe01;
			16'hdc8d: y = 16'hfe01;
			16'hdc8e: y = 16'hfe01;
			16'hdc8f: y = 16'hfe01;
			16'hdc90: y = 16'hfe01;
			16'hdc91: y = 16'hfe01;
			16'hdc92: y = 16'hfe01;
			16'hdc93: y = 16'hfe01;
			16'hdc94: y = 16'hfe01;
			16'hdc95: y = 16'hfe01;
			16'hdc96: y = 16'hfe01;
			16'hdc97: y = 16'hfe01;
			16'hdc98: y = 16'hfe01;
			16'hdc99: y = 16'hfe01;
			16'hdc9a: y = 16'hfe01;
			16'hdc9b: y = 16'hfe01;
			16'hdc9c: y = 16'hfe01;
			16'hdc9d: y = 16'hfe01;
			16'hdc9e: y = 16'hfe01;
			16'hdc9f: y = 16'hfe01;
			16'hdca0: y = 16'hfe01;
			16'hdca1: y = 16'hfe01;
			16'hdca2: y = 16'hfe01;
			16'hdca3: y = 16'hfe01;
			16'hdca4: y = 16'hfe01;
			16'hdca5: y = 16'hfe01;
			16'hdca6: y = 16'hfe01;
			16'hdca7: y = 16'hfe01;
			16'hdca8: y = 16'hfe01;
			16'hdca9: y = 16'hfe01;
			16'hdcaa: y = 16'hfe01;
			16'hdcab: y = 16'hfe01;
			16'hdcac: y = 16'hfe01;
			16'hdcad: y = 16'hfe01;
			16'hdcae: y = 16'hfe01;
			16'hdcaf: y = 16'hfe01;
			16'hdcb0: y = 16'hfe01;
			16'hdcb1: y = 16'hfe01;
			16'hdcb2: y = 16'hfe01;
			16'hdcb3: y = 16'hfe01;
			16'hdcb4: y = 16'hfe01;
			16'hdcb5: y = 16'hfe01;
			16'hdcb6: y = 16'hfe01;
			16'hdcb7: y = 16'hfe01;
			16'hdcb8: y = 16'hfe01;
			16'hdcb9: y = 16'hfe01;
			16'hdcba: y = 16'hfe01;
			16'hdcbb: y = 16'hfe01;
			16'hdcbc: y = 16'hfe01;
			16'hdcbd: y = 16'hfe01;
			16'hdcbe: y = 16'hfe01;
			16'hdcbf: y = 16'hfe01;
			16'hdcc0: y = 16'hfe01;
			16'hdcc1: y = 16'hfe01;
			16'hdcc2: y = 16'hfe01;
			16'hdcc3: y = 16'hfe01;
			16'hdcc4: y = 16'hfe01;
			16'hdcc5: y = 16'hfe01;
			16'hdcc6: y = 16'hfe01;
			16'hdcc7: y = 16'hfe01;
			16'hdcc8: y = 16'hfe01;
			16'hdcc9: y = 16'hfe01;
			16'hdcca: y = 16'hfe01;
			16'hdccb: y = 16'hfe01;
			16'hdccc: y = 16'hfe01;
			16'hdccd: y = 16'hfe01;
			16'hdcce: y = 16'hfe01;
			16'hdccf: y = 16'hfe01;
			16'hdcd0: y = 16'hfe01;
			16'hdcd1: y = 16'hfe01;
			16'hdcd2: y = 16'hfe01;
			16'hdcd3: y = 16'hfe01;
			16'hdcd4: y = 16'hfe01;
			16'hdcd5: y = 16'hfe01;
			16'hdcd6: y = 16'hfe01;
			16'hdcd7: y = 16'hfe01;
			16'hdcd8: y = 16'hfe01;
			16'hdcd9: y = 16'hfe01;
			16'hdcda: y = 16'hfe01;
			16'hdcdb: y = 16'hfe01;
			16'hdcdc: y = 16'hfe01;
			16'hdcdd: y = 16'hfe01;
			16'hdcde: y = 16'hfe01;
			16'hdcdf: y = 16'hfe01;
			16'hdce0: y = 16'hfe01;
			16'hdce1: y = 16'hfe01;
			16'hdce2: y = 16'hfe01;
			16'hdce3: y = 16'hfe01;
			16'hdce4: y = 16'hfe01;
			16'hdce5: y = 16'hfe01;
			16'hdce6: y = 16'hfe01;
			16'hdce7: y = 16'hfe01;
			16'hdce8: y = 16'hfe01;
			16'hdce9: y = 16'hfe01;
			16'hdcea: y = 16'hfe01;
			16'hdceb: y = 16'hfe01;
			16'hdcec: y = 16'hfe01;
			16'hdced: y = 16'hfe01;
			16'hdcee: y = 16'hfe01;
			16'hdcef: y = 16'hfe01;
			16'hdcf0: y = 16'hfe01;
			16'hdcf1: y = 16'hfe01;
			16'hdcf2: y = 16'hfe01;
			16'hdcf3: y = 16'hfe01;
			16'hdcf4: y = 16'hfe01;
			16'hdcf5: y = 16'hfe01;
			16'hdcf6: y = 16'hfe01;
			16'hdcf7: y = 16'hfe01;
			16'hdcf8: y = 16'hfe01;
			16'hdcf9: y = 16'hfe01;
			16'hdcfa: y = 16'hfe01;
			16'hdcfb: y = 16'hfe01;
			16'hdcfc: y = 16'hfe01;
			16'hdcfd: y = 16'hfe01;
			16'hdcfe: y = 16'hfe01;
			16'hdcff: y = 16'hfe01;
			16'hdd00: y = 16'hfe01;
			16'hdd01: y = 16'hfe01;
			16'hdd02: y = 16'hfe01;
			16'hdd03: y = 16'hfe01;
			16'hdd04: y = 16'hfe01;
			16'hdd05: y = 16'hfe01;
			16'hdd06: y = 16'hfe01;
			16'hdd07: y = 16'hfe01;
			16'hdd08: y = 16'hfe01;
			16'hdd09: y = 16'hfe01;
			16'hdd0a: y = 16'hfe01;
			16'hdd0b: y = 16'hfe01;
			16'hdd0c: y = 16'hfe01;
			16'hdd0d: y = 16'hfe01;
			16'hdd0e: y = 16'hfe01;
			16'hdd0f: y = 16'hfe01;
			16'hdd10: y = 16'hfe01;
			16'hdd11: y = 16'hfe01;
			16'hdd12: y = 16'hfe01;
			16'hdd13: y = 16'hfe01;
			16'hdd14: y = 16'hfe01;
			16'hdd15: y = 16'hfe01;
			16'hdd16: y = 16'hfe01;
			16'hdd17: y = 16'hfe01;
			16'hdd18: y = 16'hfe01;
			16'hdd19: y = 16'hfe01;
			16'hdd1a: y = 16'hfe01;
			16'hdd1b: y = 16'hfe01;
			16'hdd1c: y = 16'hfe01;
			16'hdd1d: y = 16'hfe01;
			16'hdd1e: y = 16'hfe01;
			16'hdd1f: y = 16'hfe01;
			16'hdd20: y = 16'hfe01;
			16'hdd21: y = 16'hfe01;
			16'hdd22: y = 16'hfe01;
			16'hdd23: y = 16'hfe01;
			16'hdd24: y = 16'hfe01;
			16'hdd25: y = 16'hfe01;
			16'hdd26: y = 16'hfe01;
			16'hdd27: y = 16'hfe01;
			16'hdd28: y = 16'hfe01;
			16'hdd29: y = 16'hfe01;
			16'hdd2a: y = 16'hfe01;
			16'hdd2b: y = 16'hfe01;
			16'hdd2c: y = 16'hfe01;
			16'hdd2d: y = 16'hfe01;
			16'hdd2e: y = 16'hfe01;
			16'hdd2f: y = 16'hfe01;
			16'hdd30: y = 16'hfe01;
			16'hdd31: y = 16'hfe01;
			16'hdd32: y = 16'hfe01;
			16'hdd33: y = 16'hfe01;
			16'hdd34: y = 16'hfe01;
			16'hdd35: y = 16'hfe01;
			16'hdd36: y = 16'hfe01;
			16'hdd37: y = 16'hfe01;
			16'hdd38: y = 16'hfe01;
			16'hdd39: y = 16'hfe01;
			16'hdd3a: y = 16'hfe01;
			16'hdd3b: y = 16'hfe01;
			16'hdd3c: y = 16'hfe01;
			16'hdd3d: y = 16'hfe01;
			16'hdd3e: y = 16'hfe01;
			16'hdd3f: y = 16'hfe01;
			16'hdd40: y = 16'hfe01;
			16'hdd41: y = 16'hfe01;
			16'hdd42: y = 16'hfe01;
			16'hdd43: y = 16'hfe01;
			16'hdd44: y = 16'hfe01;
			16'hdd45: y = 16'hfe01;
			16'hdd46: y = 16'hfe01;
			16'hdd47: y = 16'hfe01;
			16'hdd48: y = 16'hfe01;
			16'hdd49: y = 16'hfe01;
			16'hdd4a: y = 16'hfe01;
			16'hdd4b: y = 16'hfe01;
			16'hdd4c: y = 16'hfe01;
			16'hdd4d: y = 16'hfe01;
			16'hdd4e: y = 16'hfe01;
			16'hdd4f: y = 16'hfe01;
			16'hdd50: y = 16'hfe01;
			16'hdd51: y = 16'hfe01;
			16'hdd52: y = 16'hfe01;
			16'hdd53: y = 16'hfe01;
			16'hdd54: y = 16'hfe01;
			16'hdd55: y = 16'hfe01;
			16'hdd56: y = 16'hfe01;
			16'hdd57: y = 16'hfe01;
			16'hdd58: y = 16'hfe01;
			16'hdd59: y = 16'hfe01;
			16'hdd5a: y = 16'hfe01;
			16'hdd5b: y = 16'hfe01;
			16'hdd5c: y = 16'hfe01;
			16'hdd5d: y = 16'hfe01;
			16'hdd5e: y = 16'hfe01;
			16'hdd5f: y = 16'hfe01;
			16'hdd60: y = 16'hfe01;
			16'hdd61: y = 16'hfe01;
			16'hdd62: y = 16'hfe01;
			16'hdd63: y = 16'hfe01;
			16'hdd64: y = 16'hfe01;
			16'hdd65: y = 16'hfe01;
			16'hdd66: y = 16'hfe01;
			16'hdd67: y = 16'hfe01;
			16'hdd68: y = 16'hfe01;
			16'hdd69: y = 16'hfe01;
			16'hdd6a: y = 16'hfe01;
			16'hdd6b: y = 16'hfe01;
			16'hdd6c: y = 16'hfe01;
			16'hdd6d: y = 16'hfe01;
			16'hdd6e: y = 16'hfe01;
			16'hdd6f: y = 16'hfe01;
			16'hdd70: y = 16'hfe01;
			16'hdd71: y = 16'hfe01;
			16'hdd72: y = 16'hfe01;
			16'hdd73: y = 16'hfe01;
			16'hdd74: y = 16'hfe01;
			16'hdd75: y = 16'hfe01;
			16'hdd76: y = 16'hfe01;
			16'hdd77: y = 16'hfe01;
			16'hdd78: y = 16'hfe01;
			16'hdd79: y = 16'hfe01;
			16'hdd7a: y = 16'hfe01;
			16'hdd7b: y = 16'hfe01;
			16'hdd7c: y = 16'hfe01;
			16'hdd7d: y = 16'hfe01;
			16'hdd7e: y = 16'hfe01;
			16'hdd7f: y = 16'hfe01;
			16'hdd80: y = 16'hfe01;
			16'hdd81: y = 16'hfe01;
			16'hdd82: y = 16'hfe01;
			16'hdd83: y = 16'hfe01;
			16'hdd84: y = 16'hfe01;
			16'hdd85: y = 16'hfe01;
			16'hdd86: y = 16'hfe01;
			16'hdd87: y = 16'hfe01;
			16'hdd88: y = 16'hfe01;
			16'hdd89: y = 16'hfe01;
			16'hdd8a: y = 16'hfe01;
			16'hdd8b: y = 16'hfe01;
			16'hdd8c: y = 16'hfe01;
			16'hdd8d: y = 16'hfe01;
			16'hdd8e: y = 16'hfe01;
			16'hdd8f: y = 16'hfe01;
			16'hdd90: y = 16'hfe01;
			16'hdd91: y = 16'hfe01;
			16'hdd92: y = 16'hfe01;
			16'hdd93: y = 16'hfe01;
			16'hdd94: y = 16'hfe01;
			16'hdd95: y = 16'hfe01;
			16'hdd96: y = 16'hfe01;
			16'hdd97: y = 16'hfe01;
			16'hdd98: y = 16'hfe01;
			16'hdd99: y = 16'hfe01;
			16'hdd9a: y = 16'hfe01;
			16'hdd9b: y = 16'hfe01;
			16'hdd9c: y = 16'hfe01;
			16'hdd9d: y = 16'hfe01;
			16'hdd9e: y = 16'hfe01;
			16'hdd9f: y = 16'hfe01;
			16'hdda0: y = 16'hfe01;
			16'hdda1: y = 16'hfe01;
			16'hdda2: y = 16'hfe01;
			16'hdda3: y = 16'hfe01;
			16'hdda4: y = 16'hfe01;
			16'hdda5: y = 16'hfe01;
			16'hdda6: y = 16'hfe01;
			16'hdda7: y = 16'hfe01;
			16'hdda8: y = 16'hfe01;
			16'hdda9: y = 16'hfe01;
			16'hddaa: y = 16'hfe01;
			16'hddab: y = 16'hfe01;
			16'hddac: y = 16'hfe01;
			16'hddad: y = 16'hfe01;
			16'hddae: y = 16'hfe01;
			16'hddaf: y = 16'hfe01;
			16'hddb0: y = 16'hfe01;
			16'hddb1: y = 16'hfe01;
			16'hddb2: y = 16'hfe01;
			16'hddb3: y = 16'hfe01;
			16'hddb4: y = 16'hfe01;
			16'hddb5: y = 16'hfe01;
			16'hddb6: y = 16'hfe01;
			16'hddb7: y = 16'hfe01;
			16'hddb8: y = 16'hfe01;
			16'hddb9: y = 16'hfe01;
			16'hddba: y = 16'hfe01;
			16'hddbb: y = 16'hfe01;
			16'hddbc: y = 16'hfe01;
			16'hddbd: y = 16'hfe01;
			16'hddbe: y = 16'hfe01;
			16'hddbf: y = 16'hfe01;
			16'hddc0: y = 16'hfe01;
			16'hddc1: y = 16'hfe01;
			16'hddc2: y = 16'hfe01;
			16'hddc3: y = 16'hfe01;
			16'hddc4: y = 16'hfe01;
			16'hddc5: y = 16'hfe01;
			16'hddc6: y = 16'hfe01;
			16'hddc7: y = 16'hfe01;
			16'hddc8: y = 16'hfe01;
			16'hddc9: y = 16'hfe01;
			16'hddca: y = 16'hfe01;
			16'hddcb: y = 16'hfe01;
			16'hddcc: y = 16'hfe01;
			16'hddcd: y = 16'hfe01;
			16'hddce: y = 16'hfe01;
			16'hddcf: y = 16'hfe01;
			16'hddd0: y = 16'hfe01;
			16'hddd1: y = 16'hfe01;
			16'hddd2: y = 16'hfe01;
			16'hddd3: y = 16'hfe01;
			16'hddd4: y = 16'hfe01;
			16'hddd5: y = 16'hfe01;
			16'hddd6: y = 16'hfe01;
			16'hddd7: y = 16'hfe01;
			16'hddd8: y = 16'hfe01;
			16'hddd9: y = 16'hfe01;
			16'hddda: y = 16'hfe01;
			16'hdddb: y = 16'hfe01;
			16'hdddc: y = 16'hfe01;
			16'hdddd: y = 16'hfe01;
			16'hddde: y = 16'hfe01;
			16'hdddf: y = 16'hfe01;
			16'hdde0: y = 16'hfe01;
			16'hdde1: y = 16'hfe01;
			16'hdde2: y = 16'hfe01;
			16'hdde3: y = 16'hfe01;
			16'hdde4: y = 16'hfe01;
			16'hdde5: y = 16'hfe01;
			16'hdde6: y = 16'hfe01;
			16'hdde7: y = 16'hfe01;
			16'hdde8: y = 16'hfe01;
			16'hdde9: y = 16'hfe01;
			16'hddea: y = 16'hfe01;
			16'hddeb: y = 16'hfe01;
			16'hddec: y = 16'hfe01;
			16'hdded: y = 16'hfe01;
			16'hddee: y = 16'hfe01;
			16'hddef: y = 16'hfe01;
			16'hddf0: y = 16'hfe01;
			16'hddf1: y = 16'hfe01;
			16'hddf2: y = 16'hfe01;
			16'hddf3: y = 16'hfe01;
			16'hddf4: y = 16'hfe01;
			16'hddf5: y = 16'hfe01;
			16'hddf6: y = 16'hfe01;
			16'hddf7: y = 16'hfe01;
			16'hddf8: y = 16'hfe01;
			16'hddf9: y = 16'hfe01;
			16'hddfa: y = 16'hfe01;
			16'hddfb: y = 16'hfe01;
			16'hddfc: y = 16'hfe01;
			16'hddfd: y = 16'hfe01;
			16'hddfe: y = 16'hfe01;
			16'hddff: y = 16'hfe01;
			16'hde00: y = 16'hfe01;
			16'hde01: y = 16'hfe01;
			16'hde02: y = 16'hfe01;
			16'hde03: y = 16'hfe01;
			16'hde04: y = 16'hfe01;
			16'hde05: y = 16'hfe01;
			16'hde06: y = 16'hfe01;
			16'hde07: y = 16'hfe01;
			16'hde08: y = 16'hfe01;
			16'hde09: y = 16'hfe01;
			16'hde0a: y = 16'hfe01;
			16'hde0b: y = 16'hfe01;
			16'hde0c: y = 16'hfe01;
			16'hde0d: y = 16'hfe01;
			16'hde0e: y = 16'hfe01;
			16'hde0f: y = 16'hfe01;
			16'hde10: y = 16'hfe01;
			16'hde11: y = 16'hfe01;
			16'hde12: y = 16'hfe01;
			16'hde13: y = 16'hfe01;
			16'hde14: y = 16'hfe01;
			16'hde15: y = 16'hfe01;
			16'hde16: y = 16'hfe01;
			16'hde17: y = 16'hfe01;
			16'hde18: y = 16'hfe01;
			16'hde19: y = 16'hfe01;
			16'hde1a: y = 16'hfe01;
			16'hde1b: y = 16'hfe01;
			16'hde1c: y = 16'hfe01;
			16'hde1d: y = 16'hfe01;
			16'hde1e: y = 16'hfe01;
			16'hde1f: y = 16'hfe01;
			16'hde20: y = 16'hfe01;
			16'hde21: y = 16'hfe01;
			16'hde22: y = 16'hfe01;
			16'hde23: y = 16'hfe01;
			16'hde24: y = 16'hfe01;
			16'hde25: y = 16'hfe01;
			16'hde26: y = 16'hfe01;
			16'hde27: y = 16'hfe01;
			16'hde28: y = 16'hfe01;
			16'hde29: y = 16'hfe01;
			16'hde2a: y = 16'hfe01;
			16'hde2b: y = 16'hfe01;
			16'hde2c: y = 16'hfe01;
			16'hde2d: y = 16'hfe01;
			16'hde2e: y = 16'hfe01;
			16'hde2f: y = 16'hfe01;
			16'hde30: y = 16'hfe01;
			16'hde31: y = 16'hfe01;
			16'hde32: y = 16'hfe01;
			16'hde33: y = 16'hfe01;
			16'hde34: y = 16'hfe01;
			16'hde35: y = 16'hfe01;
			16'hde36: y = 16'hfe01;
			16'hde37: y = 16'hfe01;
			16'hde38: y = 16'hfe01;
			16'hde39: y = 16'hfe01;
			16'hde3a: y = 16'hfe01;
			16'hde3b: y = 16'hfe01;
			16'hde3c: y = 16'hfe01;
			16'hde3d: y = 16'hfe01;
			16'hde3e: y = 16'hfe01;
			16'hde3f: y = 16'hfe01;
			16'hde40: y = 16'hfe01;
			16'hde41: y = 16'hfe01;
			16'hde42: y = 16'hfe01;
			16'hde43: y = 16'hfe01;
			16'hde44: y = 16'hfe01;
			16'hde45: y = 16'hfe01;
			16'hde46: y = 16'hfe01;
			16'hde47: y = 16'hfe01;
			16'hde48: y = 16'hfe01;
			16'hde49: y = 16'hfe01;
			16'hde4a: y = 16'hfe01;
			16'hde4b: y = 16'hfe01;
			16'hde4c: y = 16'hfe01;
			16'hde4d: y = 16'hfe01;
			16'hde4e: y = 16'hfe01;
			16'hde4f: y = 16'hfe01;
			16'hde50: y = 16'hfe01;
			16'hde51: y = 16'hfe01;
			16'hde52: y = 16'hfe01;
			16'hde53: y = 16'hfe01;
			16'hde54: y = 16'hfe01;
			16'hde55: y = 16'hfe01;
			16'hde56: y = 16'hfe01;
			16'hde57: y = 16'hfe01;
			16'hde58: y = 16'hfe01;
			16'hde59: y = 16'hfe01;
			16'hde5a: y = 16'hfe01;
			16'hde5b: y = 16'hfe01;
			16'hde5c: y = 16'hfe01;
			16'hde5d: y = 16'hfe01;
			16'hde5e: y = 16'hfe01;
			16'hde5f: y = 16'hfe01;
			16'hde60: y = 16'hfe01;
			16'hde61: y = 16'hfe01;
			16'hde62: y = 16'hfe01;
			16'hde63: y = 16'hfe01;
			16'hde64: y = 16'hfe01;
			16'hde65: y = 16'hfe01;
			16'hde66: y = 16'hfe01;
			16'hde67: y = 16'hfe01;
			16'hde68: y = 16'hfe01;
			16'hde69: y = 16'hfe01;
			16'hde6a: y = 16'hfe01;
			16'hde6b: y = 16'hfe01;
			16'hde6c: y = 16'hfe01;
			16'hde6d: y = 16'hfe01;
			16'hde6e: y = 16'hfe01;
			16'hde6f: y = 16'hfe01;
			16'hde70: y = 16'hfe01;
			16'hde71: y = 16'hfe01;
			16'hde72: y = 16'hfe01;
			16'hde73: y = 16'hfe01;
			16'hde74: y = 16'hfe01;
			16'hde75: y = 16'hfe01;
			16'hde76: y = 16'hfe01;
			16'hde77: y = 16'hfe01;
			16'hde78: y = 16'hfe01;
			16'hde79: y = 16'hfe01;
			16'hde7a: y = 16'hfe01;
			16'hde7b: y = 16'hfe01;
			16'hde7c: y = 16'hfe01;
			16'hde7d: y = 16'hfe01;
			16'hde7e: y = 16'hfe01;
			16'hde7f: y = 16'hfe01;
			16'hde80: y = 16'hfe01;
			16'hde81: y = 16'hfe01;
			16'hde82: y = 16'hfe01;
			16'hde83: y = 16'hfe01;
			16'hde84: y = 16'hfe01;
			16'hde85: y = 16'hfe01;
			16'hde86: y = 16'hfe01;
			16'hde87: y = 16'hfe01;
			16'hde88: y = 16'hfe01;
			16'hde89: y = 16'hfe01;
			16'hde8a: y = 16'hfe01;
			16'hde8b: y = 16'hfe01;
			16'hde8c: y = 16'hfe01;
			16'hde8d: y = 16'hfe01;
			16'hde8e: y = 16'hfe01;
			16'hde8f: y = 16'hfe01;
			16'hde90: y = 16'hfe01;
			16'hde91: y = 16'hfe01;
			16'hde92: y = 16'hfe01;
			16'hde93: y = 16'hfe01;
			16'hde94: y = 16'hfe01;
			16'hde95: y = 16'hfe01;
			16'hde96: y = 16'hfe01;
			16'hde97: y = 16'hfe01;
			16'hde98: y = 16'hfe01;
			16'hde99: y = 16'hfe01;
			16'hde9a: y = 16'hfe01;
			16'hde9b: y = 16'hfe01;
			16'hde9c: y = 16'hfe01;
			16'hde9d: y = 16'hfe01;
			16'hde9e: y = 16'hfe01;
			16'hde9f: y = 16'hfe01;
			16'hdea0: y = 16'hfe01;
			16'hdea1: y = 16'hfe01;
			16'hdea2: y = 16'hfe01;
			16'hdea3: y = 16'hfe01;
			16'hdea4: y = 16'hfe01;
			16'hdea5: y = 16'hfe01;
			16'hdea6: y = 16'hfe01;
			16'hdea7: y = 16'hfe01;
			16'hdea8: y = 16'hfe01;
			16'hdea9: y = 16'hfe01;
			16'hdeaa: y = 16'hfe01;
			16'hdeab: y = 16'hfe01;
			16'hdeac: y = 16'hfe01;
			16'hdead: y = 16'hfe01;
			16'hdeae: y = 16'hfe01;
			16'hdeaf: y = 16'hfe01;
			16'hdeb0: y = 16'hfe01;
			16'hdeb1: y = 16'hfe01;
			16'hdeb2: y = 16'hfe01;
			16'hdeb3: y = 16'hfe01;
			16'hdeb4: y = 16'hfe01;
			16'hdeb5: y = 16'hfe01;
			16'hdeb6: y = 16'hfe01;
			16'hdeb7: y = 16'hfe01;
			16'hdeb8: y = 16'hfe01;
			16'hdeb9: y = 16'hfe01;
			16'hdeba: y = 16'hfe01;
			16'hdebb: y = 16'hfe01;
			16'hdebc: y = 16'hfe01;
			16'hdebd: y = 16'hfe01;
			16'hdebe: y = 16'hfe01;
			16'hdebf: y = 16'hfe01;
			16'hdec0: y = 16'hfe01;
			16'hdec1: y = 16'hfe01;
			16'hdec2: y = 16'hfe01;
			16'hdec3: y = 16'hfe01;
			16'hdec4: y = 16'hfe01;
			16'hdec5: y = 16'hfe01;
			16'hdec6: y = 16'hfe01;
			16'hdec7: y = 16'hfe01;
			16'hdec8: y = 16'hfe01;
			16'hdec9: y = 16'hfe01;
			16'hdeca: y = 16'hfe01;
			16'hdecb: y = 16'hfe01;
			16'hdecc: y = 16'hfe01;
			16'hdecd: y = 16'hfe01;
			16'hdece: y = 16'hfe01;
			16'hdecf: y = 16'hfe01;
			16'hded0: y = 16'hfe01;
			16'hded1: y = 16'hfe01;
			16'hded2: y = 16'hfe01;
			16'hded3: y = 16'hfe01;
			16'hded4: y = 16'hfe01;
			16'hded5: y = 16'hfe01;
			16'hded6: y = 16'hfe01;
			16'hded7: y = 16'hfe01;
			16'hded8: y = 16'hfe01;
			16'hded9: y = 16'hfe01;
			16'hdeda: y = 16'hfe01;
			16'hdedb: y = 16'hfe01;
			16'hdedc: y = 16'hfe01;
			16'hdedd: y = 16'hfe01;
			16'hdede: y = 16'hfe01;
			16'hdedf: y = 16'hfe01;
			16'hdee0: y = 16'hfe01;
			16'hdee1: y = 16'hfe01;
			16'hdee2: y = 16'hfe01;
			16'hdee3: y = 16'hfe01;
			16'hdee4: y = 16'hfe01;
			16'hdee5: y = 16'hfe01;
			16'hdee6: y = 16'hfe01;
			16'hdee7: y = 16'hfe01;
			16'hdee8: y = 16'hfe01;
			16'hdee9: y = 16'hfe01;
			16'hdeea: y = 16'hfe01;
			16'hdeeb: y = 16'hfe01;
			16'hdeec: y = 16'hfe01;
			16'hdeed: y = 16'hfe01;
			16'hdeee: y = 16'hfe01;
			16'hdeef: y = 16'hfe01;
			16'hdef0: y = 16'hfe01;
			16'hdef1: y = 16'hfe01;
			16'hdef2: y = 16'hfe01;
			16'hdef3: y = 16'hfe01;
			16'hdef4: y = 16'hfe01;
			16'hdef5: y = 16'hfe01;
			16'hdef6: y = 16'hfe01;
			16'hdef7: y = 16'hfe01;
			16'hdef8: y = 16'hfe01;
			16'hdef9: y = 16'hfe01;
			16'hdefa: y = 16'hfe01;
			16'hdefb: y = 16'hfe01;
			16'hdefc: y = 16'hfe01;
			16'hdefd: y = 16'hfe01;
			16'hdefe: y = 16'hfe01;
			16'hdeff: y = 16'hfe01;
			16'hdf00: y = 16'hfe01;
			16'hdf01: y = 16'hfe01;
			16'hdf02: y = 16'hfe01;
			16'hdf03: y = 16'hfe01;
			16'hdf04: y = 16'hfe01;
			16'hdf05: y = 16'hfe01;
			16'hdf06: y = 16'hfe01;
			16'hdf07: y = 16'hfe01;
			16'hdf08: y = 16'hfe01;
			16'hdf09: y = 16'hfe01;
			16'hdf0a: y = 16'hfe01;
			16'hdf0b: y = 16'hfe01;
			16'hdf0c: y = 16'hfe01;
			16'hdf0d: y = 16'hfe01;
			16'hdf0e: y = 16'hfe01;
			16'hdf0f: y = 16'hfe01;
			16'hdf10: y = 16'hfe01;
			16'hdf11: y = 16'hfe01;
			16'hdf12: y = 16'hfe01;
			16'hdf13: y = 16'hfe01;
			16'hdf14: y = 16'hfe01;
			16'hdf15: y = 16'hfe01;
			16'hdf16: y = 16'hfe01;
			16'hdf17: y = 16'hfe01;
			16'hdf18: y = 16'hfe01;
			16'hdf19: y = 16'hfe01;
			16'hdf1a: y = 16'hfe01;
			16'hdf1b: y = 16'hfe01;
			16'hdf1c: y = 16'hfe01;
			16'hdf1d: y = 16'hfe01;
			16'hdf1e: y = 16'hfe01;
			16'hdf1f: y = 16'hfe01;
			16'hdf20: y = 16'hfe01;
			16'hdf21: y = 16'hfe01;
			16'hdf22: y = 16'hfe01;
			16'hdf23: y = 16'hfe01;
			16'hdf24: y = 16'hfe01;
			16'hdf25: y = 16'hfe01;
			16'hdf26: y = 16'hfe01;
			16'hdf27: y = 16'hfe01;
			16'hdf28: y = 16'hfe01;
			16'hdf29: y = 16'hfe01;
			16'hdf2a: y = 16'hfe01;
			16'hdf2b: y = 16'hfe01;
			16'hdf2c: y = 16'hfe01;
			16'hdf2d: y = 16'hfe01;
			16'hdf2e: y = 16'hfe01;
			16'hdf2f: y = 16'hfe01;
			16'hdf30: y = 16'hfe01;
			16'hdf31: y = 16'hfe01;
			16'hdf32: y = 16'hfe01;
			16'hdf33: y = 16'hfe01;
			16'hdf34: y = 16'hfe01;
			16'hdf35: y = 16'hfe01;
			16'hdf36: y = 16'hfe01;
			16'hdf37: y = 16'hfe01;
			16'hdf38: y = 16'hfe01;
			16'hdf39: y = 16'hfe01;
			16'hdf3a: y = 16'hfe01;
			16'hdf3b: y = 16'hfe01;
			16'hdf3c: y = 16'hfe01;
			16'hdf3d: y = 16'hfe01;
			16'hdf3e: y = 16'hfe01;
			16'hdf3f: y = 16'hfe01;
			16'hdf40: y = 16'hfe01;
			16'hdf41: y = 16'hfe01;
			16'hdf42: y = 16'hfe01;
			16'hdf43: y = 16'hfe01;
			16'hdf44: y = 16'hfe01;
			16'hdf45: y = 16'hfe01;
			16'hdf46: y = 16'hfe01;
			16'hdf47: y = 16'hfe01;
			16'hdf48: y = 16'hfe01;
			16'hdf49: y = 16'hfe01;
			16'hdf4a: y = 16'hfe01;
			16'hdf4b: y = 16'hfe01;
			16'hdf4c: y = 16'hfe01;
			16'hdf4d: y = 16'hfe01;
			16'hdf4e: y = 16'hfe01;
			16'hdf4f: y = 16'hfe01;
			16'hdf50: y = 16'hfe01;
			16'hdf51: y = 16'hfe01;
			16'hdf52: y = 16'hfe01;
			16'hdf53: y = 16'hfe01;
			16'hdf54: y = 16'hfe01;
			16'hdf55: y = 16'hfe01;
			16'hdf56: y = 16'hfe01;
			16'hdf57: y = 16'hfe01;
			16'hdf58: y = 16'hfe01;
			16'hdf59: y = 16'hfe01;
			16'hdf5a: y = 16'hfe01;
			16'hdf5b: y = 16'hfe01;
			16'hdf5c: y = 16'hfe01;
			16'hdf5d: y = 16'hfe01;
			16'hdf5e: y = 16'hfe01;
			16'hdf5f: y = 16'hfe01;
			16'hdf60: y = 16'hfe01;
			16'hdf61: y = 16'hfe01;
			16'hdf62: y = 16'hfe01;
			16'hdf63: y = 16'hfe01;
			16'hdf64: y = 16'hfe01;
			16'hdf65: y = 16'hfe01;
			16'hdf66: y = 16'hfe01;
			16'hdf67: y = 16'hfe01;
			16'hdf68: y = 16'hfe01;
			16'hdf69: y = 16'hfe01;
			16'hdf6a: y = 16'hfe01;
			16'hdf6b: y = 16'hfe01;
			16'hdf6c: y = 16'hfe01;
			16'hdf6d: y = 16'hfe01;
			16'hdf6e: y = 16'hfe01;
			16'hdf6f: y = 16'hfe01;
			16'hdf70: y = 16'hfe01;
			16'hdf71: y = 16'hfe01;
			16'hdf72: y = 16'hfe01;
			16'hdf73: y = 16'hfe01;
			16'hdf74: y = 16'hfe01;
			16'hdf75: y = 16'hfe01;
			16'hdf76: y = 16'hfe01;
			16'hdf77: y = 16'hfe01;
			16'hdf78: y = 16'hfe01;
			16'hdf79: y = 16'hfe01;
			16'hdf7a: y = 16'hfe01;
			16'hdf7b: y = 16'hfe01;
			16'hdf7c: y = 16'hfe01;
			16'hdf7d: y = 16'hfe01;
			16'hdf7e: y = 16'hfe01;
			16'hdf7f: y = 16'hfe01;
			16'hdf80: y = 16'hfe01;
			16'hdf81: y = 16'hfe01;
			16'hdf82: y = 16'hfe01;
			16'hdf83: y = 16'hfe01;
			16'hdf84: y = 16'hfe01;
			16'hdf85: y = 16'hfe01;
			16'hdf86: y = 16'hfe01;
			16'hdf87: y = 16'hfe01;
			16'hdf88: y = 16'hfe01;
			16'hdf89: y = 16'hfe01;
			16'hdf8a: y = 16'hfe01;
			16'hdf8b: y = 16'hfe01;
			16'hdf8c: y = 16'hfe01;
			16'hdf8d: y = 16'hfe01;
			16'hdf8e: y = 16'hfe01;
			16'hdf8f: y = 16'hfe01;
			16'hdf90: y = 16'hfe01;
			16'hdf91: y = 16'hfe01;
			16'hdf92: y = 16'hfe01;
			16'hdf93: y = 16'hfe01;
			16'hdf94: y = 16'hfe01;
			16'hdf95: y = 16'hfe01;
			16'hdf96: y = 16'hfe01;
			16'hdf97: y = 16'hfe01;
			16'hdf98: y = 16'hfe01;
			16'hdf99: y = 16'hfe01;
			16'hdf9a: y = 16'hfe01;
			16'hdf9b: y = 16'hfe01;
			16'hdf9c: y = 16'hfe01;
			16'hdf9d: y = 16'hfe01;
			16'hdf9e: y = 16'hfe01;
			16'hdf9f: y = 16'hfe01;
			16'hdfa0: y = 16'hfe01;
			16'hdfa1: y = 16'hfe01;
			16'hdfa2: y = 16'hfe01;
			16'hdfa3: y = 16'hfe01;
			16'hdfa4: y = 16'hfe01;
			16'hdfa5: y = 16'hfe01;
			16'hdfa6: y = 16'hfe01;
			16'hdfa7: y = 16'hfe01;
			16'hdfa8: y = 16'hfe01;
			16'hdfa9: y = 16'hfe01;
			16'hdfaa: y = 16'hfe01;
			16'hdfab: y = 16'hfe01;
			16'hdfac: y = 16'hfe01;
			16'hdfad: y = 16'hfe01;
			16'hdfae: y = 16'hfe01;
			16'hdfaf: y = 16'hfe01;
			16'hdfb0: y = 16'hfe01;
			16'hdfb1: y = 16'hfe01;
			16'hdfb2: y = 16'hfe01;
			16'hdfb3: y = 16'hfe01;
			16'hdfb4: y = 16'hfe01;
			16'hdfb5: y = 16'hfe01;
			16'hdfb6: y = 16'hfe01;
			16'hdfb7: y = 16'hfe01;
			16'hdfb8: y = 16'hfe01;
			16'hdfb9: y = 16'hfe01;
			16'hdfba: y = 16'hfe01;
			16'hdfbb: y = 16'hfe01;
			16'hdfbc: y = 16'hfe01;
			16'hdfbd: y = 16'hfe01;
			16'hdfbe: y = 16'hfe01;
			16'hdfbf: y = 16'hfe01;
			16'hdfc0: y = 16'hfe01;
			16'hdfc1: y = 16'hfe01;
			16'hdfc2: y = 16'hfe01;
			16'hdfc3: y = 16'hfe01;
			16'hdfc4: y = 16'hfe01;
			16'hdfc5: y = 16'hfe01;
			16'hdfc6: y = 16'hfe01;
			16'hdfc7: y = 16'hfe01;
			16'hdfc8: y = 16'hfe01;
			16'hdfc9: y = 16'hfe01;
			16'hdfca: y = 16'hfe01;
			16'hdfcb: y = 16'hfe01;
			16'hdfcc: y = 16'hfe01;
			16'hdfcd: y = 16'hfe01;
			16'hdfce: y = 16'hfe01;
			16'hdfcf: y = 16'hfe01;
			16'hdfd0: y = 16'hfe01;
			16'hdfd1: y = 16'hfe01;
			16'hdfd2: y = 16'hfe01;
			16'hdfd3: y = 16'hfe01;
			16'hdfd4: y = 16'hfe01;
			16'hdfd5: y = 16'hfe01;
			16'hdfd6: y = 16'hfe01;
			16'hdfd7: y = 16'hfe01;
			16'hdfd8: y = 16'hfe01;
			16'hdfd9: y = 16'hfe01;
			16'hdfda: y = 16'hfe01;
			16'hdfdb: y = 16'hfe01;
			16'hdfdc: y = 16'hfe01;
			16'hdfdd: y = 16'hfe01;
			16'hdfde: y = 16'hfe01;
			16'hdfdf: y = 16'hfe01;
			16'hdfe0: y = 16'hfe01;
			16'hdfe1: y = 16'hfe01;
			16'hdfe2: y = 16'hfe01;
			16'hdfe3: y = 16'hfe01;
			16'hdfe4: y = 16'hfe01;
			16'hdfe5: y = 16'hfe01;
			16'hdfe6: y = 16'hfe01;
			16'hdfe7: y = 16'hfe01;
			16'hdfe8: y = 16'hfe01;
			16'hdfe9: y = 16'hfe01;
			16'hdfea: y = 16'hfe01;
			16'hdfeb: y = 16'hfe01;
			16'hdfec: y = 16'hfe01;
			16'hdfed: y = 16'hfe01;
			16'hdfee: y = 16'hfe01;
			16'hdfef: y = 16'hfe01;
			16'hdff0: y = 16'hfe01;
			16'hdff1: y = 16'hfe01;
			16'hdff2: y = 16'hfe01;
			16'hdff3: y = 16'hfe01;
			16'hdff4: y = 16'hfe01;
			16'hdff5: y = 16'hfe01;
			16'hdff6: y = 16'hfe01;
			16'hdff7: y = 16'hfe01;
			16'hdff8: y = 16'hfe01;
			16'hdff9: y = 16'hfe01;
			16'hdffa: y = 16'hfe01;
			16'hdffb: y = 16'hfe01;
			16'hdffc: y = 16'hfe01;
			16'hdffd: y = 16'hfe01;
			16'hdffe: y = 16'hfe01;
			16'hdfff: y = 16'hfe01;
			16'he000: y = 16'hfe01;
			16'he001: y = 16'hfe01;
			16'he002: y = 16'hfe01;
			16'he003: y = 16'hfe01;
			16'he004: y = 16'hfe01;
			16'he005: y = 16'hfe01;
			16'he006: y = 16'hfe01;
			16'he007: y = 16'hfe01;
			16'he008: y = 16'hfe01;
			16'he009: y = 16'hfe01;
			16'he00a: y = 16'hfe01;
			16'he00b: y = 16'hfe01;
			16'he00c: y = 16'hfe01;
			16'he00d: y = 16'hfe01;
			16'he00e: y = 16'hfe01;
			16'he00f: y = 16'hfe01;
			16'he010: y = 16'hfe01;
			16'he011: y = 16'hfe01;
			16'he012: y = 16'hfe01;
			16'he013: y = 16'hfe01;
			16'he014: y = 16'hfe01;
			16'he015: y = 16'hfe01;
			16'he016: y = 16'hfe01;
			16'he017: y = 16'hfe01;
			16'he018: y = 16'hfe01;
			16'he019: y = 16'hfe01;
			16'he01a: y = 16'hfe01;
			16'he01b: y = 16'hfe01;
			16'he01c: y = 16'hfe01;
			16'he01d: y = 16'hfe01;
			16'he01e: y = 16'hfe01;
			16'he01f: y = 16'hfe01;
			16'he020: y = 16'hfe01;
			16'he021: y = 16'hfe01;
			16'he022: y = 16'hfe01;
			16'he023: y = 16'hfe01;
			16'he024: y = 16'hfe01;
			16'he025: y = 16'hfe01;
			16'he026: y = 16'hfe01;
			16'he027: y = 16'hfe01;
			16'he028: y = 16'hfe01;
			16'he029: y = 16'hfe01;
			16'he02a: y = 16'hfe01;
			16'he02b: y = 16'hfe01;
			16'he02c: y = 16'hfe01;
			16'he02d: y = 16'hfe01;
			16'he02e: y = 16'hfe01;
			16'he02f: y = 16'hfe01;
			16'he030: y = 16'hfe01;
			16'he031: y = 16'hfe01;
			16'he032: y = 16'hfe01;
			16'he033: y = 16'hfe01;
			16'he034: y = 16'hfe01;
			16'he035: y = 16'hfe01;
			16'he036: y = 16'hfe01;
			16'he037: y = 16'hfe01;
			16'he038: y = 16'hfe01;
			16'he039: y = 16'hfe01;
			16'he03a: y = 16'hfe01;
			16'he03b: y = 16'hfe01;
			16'he03c: y = 16'hfe01;
			16'he03d: y = 16'hfe01;
			16'he03e: y = 16'hfe01;
			16'he03f: y = 16'hfe01;
			16'he040: y = 16'hfe01;
			16'he041: y = 16'hfe01;
			16'he042: y = 16'hfe01;
			16'he043: y = 16'hfe01;
			16'he044: y = 16'hfe01;
			16'he045: y = 16'hfe01;
			16'he046: y = 16'hfe01;
			16'he047: y = 16'hfe01;
			16'he048: y = 16'hfe01;
			16'he049: y = 16'hfe01;
			16'he04a: y = 16'hfe01;
			16'he04b: y = 16'hfe01;
			16'he04c: y = 16'hfe01;
			16'he04d: y = 16'hfe01;
			16'he04e: y = 16'hfe01;
			16'he04f: y = 16'hfe01;
			16'he050: y = 16'hfe01;
			16'he051: y = 16'hfe01;
			16'he052: y = 16'hfe01;
			16'he053: y = 16'hfe01;
			16'he054: y = 16'hfe01;
			16'he055: y = 16'hfe01;
			16'he056: y = 16'hfe01;
			16'he057: y = 16'hfe01;
			16'he058: y = 16'hfe01;
			16'he059: y = 16'hfe01;
			16'he05a: y = 16'hfe01;
			16'he05b: y = 16'hfe01;
			16'he05c: y = 16'hfe01;
			16'he05d: y = 16'hfe01;
			16'he05e: y = 16'hfe01;
			16'he05f: y = 16'hfe01;
			16'he060: y = 16'hfe01;
			16'he061: y = 16'hfe01;
			16'he062: y = 16'hfe01;
			16'he063: y = 16'hfe01;
			16'he064: y = 16'hfe01;
			16'he065: y = 16'hfe01;
			16'he066: y = 16'hfe01;
			16'he067: y = 16'hfe01;
			16'he068: y = 16'hfe01;
			16'he069: y = 16'hfe01;
			16'he06a: y = 16'hfe01;
			16'he06b: y = 16'hfe01;
			16'he06c: y = 16'hfe01;
			16'he06d: y = 16'hfe01;
			16'he06e: y = 16'hfe01;
			16'he06f: y = 16'hfe01;
			16'he070: y = 16'hfe01;
			16'he071: y = 16'hfe01;
			16'he072: y = 16'hfe01;
			16'he073: y = 16'hfe01;
			16'he074: y = 16'hfe01;
			16'he075: y = 16'hfe01;
			16'he076: y = 16'hfe01;
			16'he077: y = 16'hfe01;
			16'he078: y = 16'hfe01;
			16'he079: y = 16'hfe01;
			16'he07a: y = 16'hfe01;
			16'he07b: y = 16'hfe01;
			16'he07c: y = 16'hfe01;
			16'he07d: y = 16'hfe01;
			16'he07e: y = 16'hfe01;
			16'he07f: y = 16'hfe01;
			16'he080: y = 16'hfe01;
			16'he081: y = 16'hfe01;
			16'he082: y = 16'hfe01;
			16'he083: y = 16'hfe01;
			16'he084: y = 16'hfe01;
			16'he085: y = 16'hfe01;
			16'he086: y = 16'hfe01;
			16'he087: y = 16'hfe01;
			16'he088: y = 16'hfe01;
			16'he089: y = 16'hfe01;
			16'he08a: y = 16'hfe01;
			16'he08b: y = 16'hfe01;
			16'he08c: y = 16'hfe01;
			16'he08d: y = 16'hfe01;
			16'he08e: y = 16'hfe01;
			16'he08f: y = 16'hfe01;
			16'he090: y = 16'hfe01;
			16'he091: y = 16'hfe01;
			16'he092: y = 16'hfe01;
			16'he093: y = 16'hfe01;
			16'he094: y = 16'hfe01;
			16'he095: y = 16'hfe01;
			16'he096: y = 16'hfe01;
			16'he097: y = 16'hfe01;
			16'he098: y = 16'hfe01;
			16'he099: y = 16'hfe01;
			16'he09a: y = 16'hfe01;
			16'he09b: y = 16'hfe01;
			16'he09c: y = 16'hfe01;
			16'he09d: y = 16'hfe01;
			16'he09e: y = 16'hfe01;
			16'he09f: y = 16'hfe01;
			16'he0a0: y = 16'hfe01;
			16'he0a1: y = 16'hfe01;
			16'he0a2: y = 16'hfe01;
			16'he0a3: y = 16'hfe01;
			16'he0a4: y = 16'hfe01;
			16'he0a5: y = 16'hfe01;
			16'he0a6: y = 16'hfe01;
			16'he0a7: y = 16'hfe01;
			16'he0a8: y = 16'hfe01;
			16'he0a9: y = 16'hfe01;
			16'he0aa: y = 16'hfe01;
			16'he0ab: y = 16'hfe01;
			16'he0ac: y = 16'hfe01;
			16'he0ad: y = 16'hfe01;
			16'he0ae: y = 16'hfe01;
			16'he0af: y = 16'hfe01;
			16'he0b0: y = 16'hfe01;
			16'he0b1: y = 16'hfe01;
			16'he0b2: y = 16'hfe01;
			16'he0b3: y = 16'hfe01;
			16'he0b4: y = 16'hfe01;
			16'he0b5: y = 16'hfe01;
			16'he0b6: y = 16'hfe01;
			16'he0b7: y = 16'hfe01;
			16'he0b8: y = 16'hfe01;
			16'he0b9: y = 16'hfe01;
			16'he0ba: y = 16'hfe01;
			16'he0bb: y = 16'hfe01;
			16'he0bc: y = 16'hfe01;
			16'he0bd: y = 16'hfe01;
			16'he0be: y = 16'hfe01;
			16'he0bf: y = 16'hfe01;
			16'he0c0: y = 16'hfe01;
			16'he0c1: y = 16'hfe01;
			16'he0c2: y = 16'hfe01;
			16'he0c3: y = 16'hfe01;
			16'he0c4: y = 16'hfe01;
			16'he0c5: y = 16'hfe01;
			16'he0c6: y = 16'hfe01;
			16'he0c7: y = 16'hfe01;
			16'he0c8: y = 16'hfe01;
			16'he0c9: y = 16'hfe01;
			16'he0ca: y = 16'hfe01;
			16'he0cb: y = 16'hfe01;
			16'he0cc: y = 16'hfe01;
			16'he0cd: y = 16'hfe01;
			16'he0ce: y = 16'hfe01;
			16'he0cf: y = 16'hfe01;
			16'he0d0: y = 16'hfe01;
			16'he0d1: y = 16'hfe01;
			16'he0d2: y = 16'hfe01;
			16'he0d3: y = 16'hfe01;
			16'he0d4: y = 16'hfe01;
			16'he0d5: y = 16'hfe01;
			16'he0d6: y = 16'hfe01;
			16'he0d7: y = 16'hfe01;
			16'he0d8: y = 16'hfe01;
			16'he0d9: y = 16'hfe01;
			16'he0da: y = 16'hfe01;
			16'he0db: y = 16'hfe01;
			16'he0dc: y = 16'hfe01;
			16'he0dd: y = 16'hfe01;
			16'he0de: y = 16'hfe01;
			16'he0df: y = 16'hfe01;
			16'he0e0: y = 16'hfe01;
			16'he0e1: y = 16'hfe01;
			16'he0e2: y = 16'hfe01;
			16'he0e3: y = 16'hfe01;
			16'he0e4: y = 16'hfe01;
			16'he0e5: y = 16'hfe01;
			16'he0e6: y = 16'hfe01;
			16'he0e7: y = 16'hfe01;
			16'he0e8: y = 16'hfe01;
			16'he0e9: y = 16'hfe01;
			16'he0ea: y = 16'hfe01;
			16'he0eb: y = 16'hfe01;
			16'he0ec: y = 16'hfe01;
			16'he0ed: y = 16'hfe01;
			16'he0ee: y = 16'hfe01;
			16'he0ef: y = 16'hfe01;
			16'he0f0: y = 16'hfe01;
			16'he0f1: y = 16'hfe01;
			16'he0f2: y = 16'hfe01;
			16'he0f3: y = 16'hfe01;
			16'he0f4: y = 16'hfe01;
			16'he0f5: y = 16'hfe01;
			16'he0f6: y = 16'hfe01;
			16'he0f7: y = 16'hfe01;
			16'he0f8: y = 16'hfe01;
			16'he0f9: y = 16'hfe01;
			16'he0fa: y = 16'hfe01;
			16'he0fb: y = 16'hfe01;
			16'he0fc: y = 16'hfe01;
			16'he0fd: y = 16'hfe01;
			16'he0fe: y = 16'hfe01;
			16'he0ff: y = 16'hfe01;
			16'he100: y = 16'hfe01;
			16'he101: y = 16'hfe01;
			16'he102: y = 16'hfe01;
			16'he103: y = 16'hfe01;
			16'he104: y = 16'hfe01;
			16'he105: y = 16'hfe01;
			16'he106: y = 16'hfe01;
			16'he107: y = 16'hfe01;
			16'he108: y = 16'hfe01;
			16'he109: y = 16'hfe01;
			16'he10a: y = 16'hfe01;
			16'he10b: y = 16'hfe01;
			16'he10c: y = 16'hfe01;
			16'he10d: y = 16'hfe01;
			16'he10e: y = 16'hfe01;
			16'he10f: y = 16'hfe01;
			16'he110: y = 16'hfe01;
			16'he111: y = 16'hfe01;
			16'he112: y = 16'hfe01;
			16'he113: y = 16'hfe01;
			16'he114: y = 16'hfe01;
			16'he115: y = 16'hfe01;
			16'he116: y = 16'hfe01;
			16'he117: y = 16'hfe01;
			16'he118: y = 16'hfe01;
			16'he119: y = 16'hfe01;
			16'he11a: y = 16'hfe01;
			16'he11b: y = 16'hfe01;
			16'he11c: y = 16'hfe01;
			16'he11d: y = 16'hfe01;
			16'he11e: y = 16'hfe01;
			16'he11f: y = 16'hfe01;
			16'he120: y = 16'hfe01;
			16'he121: y = 16'hfe01;
			16'he122: y = 16'hfe01;
			16'he123: y = 16'hfe01;
			16'he124: y = 16'hfe01;
			16'he125: y = 16'hfe01;
			16'he126: y = 16'hfe01;
			16'he127: y = 16'hfe01;
			16'he128: y = 16'hfe01;
			16'he129: y = 16'hfe01;
			16'he12a: y = 16'hfe01;
			16'he12b: y = 16'hfe01;
			16'he12c: y = 16'hfe01;
			16'he12d: y = 16'hfe01;
			16'he12e: y = 16'hfe01;
			16'he12f: y = 16'hfe01;
			16'he130: y = 16'hfe01;
			16'he131: y = 16'hfe01;
			16'he132: y = 16'hfe01;
			16'he133: y = 16'hfe01;
			16'he134: y = 16'hfe01;
			16'he135: y = 16'hfe01;
			16'he136: y = 16'hfe01;
			16'he137: y = 16'hfe01;
			16'he138: y = 16'hfe01;
			16'he139: y = 16'hfe01;
			16'he13a: y = 16'hfe01;
			16'he13b: y = 16'hfe01;
			16'he13c: y = 16'hfe01;
			16'he13d: y = 16'hfe01;
			16'he13e: y = 16'hfe01;
			16'he13f: y = 16'hfe01;
			16'he140: y = 16'hfe01;
			16'he141: y = 16'hfe01;
			16'he142: y = 16'hfe01;
			16'he143: y = 16'hfe01;
			16'he144: y = 16'hfe01;
			16'he145: y = 16'hfe01;
			16'he146: y = 16'hfe01;
			16'he147: y = 16'hfe01;
			16'he148: y = 16'hfe01;
			16'he149: y = 16'hfe01;
			16'he14a: y = 16'hfe01;
			16'he14b: y = 16'hfe01;
			16'he14c: y = 16'hfe01;
			16'he14d: y = 16'hfe01;
			16'he14e: y = 16'hfe01;
			16'he14f: y = 16'hfe01;
			16'he150: y = 16'hfe01;
			16'he151: y = 16'hfe01;
			16'he152: y = 16'hfe01;
			16'he153: y = 16'hfe01;
			16'he154: y = 16'hfe01;
			16'he155: y = 16'hfe01;
			16'he156: y = 16'hfe01;
			16'he157: y = 16'hfe01;
			16'he158: y = 16'hfe01;
			16'he159: y = 16'hfe01;
			16'he15a: y = 16'hfe01;
			16'he15b: y = 16'hfe01;
			16'he15c: y = 16'hfe01;
			16'he15d: y = 16'hfe01;
			16'he15e: y = 16'hfe01;
			16'he15f: y = 16'hfe01;
			16'he160: y = 16'hfe01;
			16'he161: y = 16'hfe01;
			16'he162: y = 16'hfe01;
			16'he163: y = 16'hfe01;
			16'he164: y = 16'hfe01;
			16'he165: y = 16'hfe01;
			16'he166: y = 16'hfe01;
			16'he167: y = 16'hfe01;
			16'he168: y = 16'hfe01;
			16'he169: y = 16'hfe01;
			16'he16a: y = 16'hfe01;
			16'he16b: y = 16'hfe01;
			16'he16c: y = 16'hfe01;
			16'he16d: y = 16'hfe01;
			16'he16e: y = 16'hfe01;
			16'he16f: y = 16'hfe01;
			16'he170: y = 16'hfe01;
			16'he171: y = 16'hfe01;
			16'he172: y = 16'hfe01;
			16'he173: y = 16'hfe01;
			16'he174: y = 16'hfe01;
			16'he175: y = 16'hfe01;
			16'he176: y = 16'hfe01;
			16'he177: y = 16'hfe01;
			16'he178: y = 16'hfe01;
			16'he179: y = 16'hfe01;
			16'he17a: y = 16'hfe01;
			16'he17b: y = 16'hfe01;
			16'he17c: y = 16'hfe01;
			16'he17d: y = 16'hfe01;
			16'he17e: y = 16'hfe01;
			16'he17f: y = 16'hfe01;
			16'he180: y = 16'hfe01;
			16'he181: y = 16'hfe01;
			16'he182: y = 16'hfe01;
			16'he183: y = 16'hfe01;
			16'he184: y = 16'hfe01;
			16'he185: y = 16'hfe01;
			16'he186: y = 16'hfe01;
			16'he187: y = 16'hfe01;
			16'he188: y = 16'hfe01;
			16'he189: y = 16'hfe01;
			16'he18a: y = 16'hfe01;
			16'he18b: y = 16'hfe01;
			16'he18c: y = 16'hfe01;
			16'he18d: y = 16'hfe01;
			16'he18e: y = 16'hfe01;
			16'he18f: y = 16'hfe01;
			16'he190: y = 16'hfe01;
			16'he191: y = 16'hfe01;
			16'he192: y = 16'hfe01;
			16'he193: y = 16'hfe01;
			16'he194: y = 16'hfe01;
			16'he195: y = 16'hfe01;
			16'he196: y = 16'hfe01;
			16'he197: y = 16'hfe01;
			16'he198: y = 16'hfe01;
			16'he199: y = 16'hfe01;
			16'he19a: y = 16'hfe01;
			16'he19b: y = 16'hfe01;
			16'he19c: y = 16'hfe01;
			16'he19d: y = 16'hfe01;
			16'he19e: y = 16'hfe01;
			16'he19f: y = 16'hfe01;
			16'he1a0: y = 16'hfe01;
			16'he1a1: y = 16'hfe01;
			16'he1a2: y = 16'hfe01;
			16'he1a3: y = 16'hfe01;
			16'he1a4: y = 16'hfe01;
			16'he1a5: y = 16'hfe01;
			16'he1a6: y = 16'hfe01;
			16'he1a7: y = 16'hfe01;
			16'he1a8: y = 16'hfe01;
			16'he1a9: y = 16'hfe01;
			16'he1aa: y = 16'hfe01;
			16'he1ab: y = 16'hfe01;
			16'he1ac: y = 16'hfe01;
			16'he1ad: y = 16'hfe01;
			16'he1ae: y = 16'hfe01;
			16'he1af: y = 16'hfe01;
			16'he1b0: y = 16'hfe01;
			16'he1b1: y = 16'hfe01;
			16'he1b2: y = 16'hfe01;
			16'he1b3: y = 16'hfe01;
			16'he1b4: y = 16'hfe01;
			16'he1b5: y = 16'hfe01;
			16'he1b6: y = 16'hfe01;
			16'he1b7: y = 16'hfe01;
			16'he1b8: y = 16'hfe01;
			16'he1b9: y = 16'hfe01;
			16'he1ba: y = 16'hfe01;
			16'he1bb: y = 16'hfe01;
			16'he1bc: y = 16'hfe01;
			16'he1bd: y = 16'hfe01;
			16'he1be: y = 16'hfe01;
			16'he1bf: y = 16'hfe01;
			16'he1c0: y = 16'hfe01;
			16'he1c1: y = 16'hfe01;
			16'he1c2: y = 16'hfe01;
			16'he1c3: y = 16'hfe01;
			16'he1c4: y = 16'hfe01;
			16'he1c5: y = 16'hfe01;
			16'he1c6: y = 16'hfe01;
			16'he1c7: y = 16'hfe01;
			16'he1c8: y = 16'hfe01;
			16'he1c9: y = 16'hfe01;
			16'he1ca: y = 16'hfe01;
			16'he1cb: y = 16'hfe01;
			16'he1cc: y = 16'hfe01;
			16'he1cd: y = 16'hfe01;
			16'he1ce: y = 16'hfe01;
			16'he1cf: y = 16'hfe01;
			16'he1d0: y = 16'hfe01;
			16'he1d1: y = 16'hfe01;
			16'he1d2: y = 16'hfe01;
			16'he1d3: y = 16'hfe01;
			16'he1d4: y = 16'hfe01;
			16'he1d5: y = 16'hfe01;
			16'he1d6: y = 16'hfe01;
			16'he1d7: y = 16'hfe01;
			16'he1d8: y = 16'hfe01;
			16'he1d9: y = 16'hfe01;
			16'he1da: y = 16'hfe01;
			16'he1db: y = 16'hfe01;
			16'he1dc: y = 16'hfe01;
			16'he1dd: y = 16'hfe01;
			16'he1de: y = 16'hfe01;
			16'he1df: y = 16'hfe01;
			16'he1e0: y = 16'hfe01;
			16'he1e1: y = 16'hfe01;
			16'he1e2: y = 16'hfe01;
			16'he1e3: y = 16'hfe01;
			16'he1e4: y = 16'hfe01;
			16'he1e5: y = 16'hfe01;
			16'he1e6: y = 16'hfe01;
			16'he1e7: y = 16'hfe01;
			16'he1e8: y = 16'hfe01;
			16'he1e9: y = 16'hfe01;
			16'he1ea: y = 16'hfe01;
			16'he1eb: y = 16'hfe01;
			16'he1ec: y = 16'hfe01;
			16'he1ed: y = 16'hfe01;
			16'he1ee: y = 16'hfe01;
			16'he1ef: y = 16'hfe01;
			16'he1f0: y = 16'hfe01;
			16'he1f1: y = 16'hfe01;
			16'he1f2: y = 16'hfe01;
			16'he1f3: y = 16'hfe01;
			16'he1f4: y = 16'hfe01;
			16'he1f5: y = 16'hfe01;
			16'he1f6: y = 16'hfe01;
			16'he1f7: y = 16'hfe01;
			16'he1f8: y = 16'hfe01;
			16'he1f9: y = 16'hfe01;
			16'he1fa: y = 16'hfe01;
			16'he1fb: y = 16'hfe01;
			16'he1fc: y = 16'hfe01;
			16'he1fd: y = 16'hfe01;
			16'he1fe: y = 16'hfe01;
			16'he1ff: y = 16'hfe01;
			16'he200: y = 16'hfe01;
			16'he201: y = 16'hfe01;
			16'he202: y = 16'hfe01;
			16'he203: y = 16'hfe01;
			16'he204: y = 16'hfe01;
			16'he205: y = 16'hfe01;
			16'he206: y = 16'hfe01;
			16'he207: y = 16'hfe01;
			16'he208: y = 16'hfe01;
			16'he209: y = 16'hfe01;
			16'he20a: y = 16'hfe01;
			16'he20b: y = 16'hfe01;
			16'he20c: y = 16'hfe01;
			16'he20d: y = 16'hfe01;
			16'he20e: y = 16'hfe01;
			16'he20f: y = 16'hfe01;
			16'he210: y = 16'hfe01;
			16'he211: y = 16'hfe01;
			16'he212: y = 16'hfe01;
			16'he213: y = 16'hfe01;
			16'he214: y = 16'hfe01;
			16'he215: y = 16'hfe01;
			16'he216: y = 16'hfe01;
			16'he217: y = 16'hfe01;
			16'he218: y = 16'hfe01;
			16'he219: y = 16'hfe01;
			16'he21a: y = 16'hfe01;
			16'he21b: y = 16'hfe01;
			16'he21c: y = 16'hfe01;
			16'he21d: y = 16'hfe01;
			16'he21e: y = 16'hfe01;
			16'he21f: y = 16'hfe01;
			16'he220: y = 16'hfe01;
			16'he221: y = 16'hfe01;
			16'he222: y = 16'hfe01;
			16'he223: y = 16'hfe01;
			16'he224: y = 16'hfe01;
			16'he225: y = 16'hfe01;
			16'he226: y = 16'hfe01;
			16'he227: y = 16'hfe01;
			16'he228: y = 16'hfe01;
			16'he229: y = 16'hfe01;
			16'he22a: y = 16'hfe01;
			16'he22b: y = 16'hfe01;
			16'he22c: y = 16'hfe01;
			16'he22d: y = 16'hfe01;
			16'he22e: y = 16'hfe01;
			16'he22f: y = 16'hfe01;
			16'he230: y = 16'hfe01;
			16'he231: y = 16'hfe01;
			16'he232: y = 16'hfe01;
			16'he233: y = 16'hfe01;
			16'he234: y = 16'hfe01;
			16'he235: y = 16'hfe01;
			16'he236: y = 16'hfe01;
			16'he237: y = 16'hfe01;
			16'he238: y = 16'hfe01;
			16'he239: y = 16'hfe01;
			16'he23a: y = 16'hfe01;
			16'he23b: y = 16'hfe01;
			16'he23c: y = 16'hfe01;
			16'he23d: y = 16'hfe01;
			16'he23e: y = 16'hfe01;
			16'he23f: y = 16'hfe01;
			16'he240: y = 16'hfe01;
			16'he241: y = 16'hfe01;
			16'he242: y = 16'hfe01;
			16'he243: y = 16'hfe01;
			16'he244: y = 16'hfe01;
			16'he245: y = 16'hfe01;
			16'he246: y = 16'hfe01;
			16'he247: y = 16'hfe01;
			16'he248: y = 16'hfe01;
			16'he249: y = 16'hfe01;
			16'he24a: y = 16'hfe01;
			16'he24b: y = 16'hfe01;
			16'he24c: y = 16'hfe01;
			16'he24d: y = 16'hfe01;
			16'he24e: y = 16'hfe01;
			16'he24f: y = 16'hfe01;
			16'he250: y = 16'hfe01;
			16'he251: y = 16'hfe01;
			16'he252: y = 16'hfe01;
			16'he253: y = 16'hfe01;
			16'he254: y = 16'hfe01;
			16'he255: y = 16'hfe01;
			16'he256: y = 16'hfe01;
			16'he257: y = 16'hfe01;
			16'he258: y = 16'hfe01;
			16'he259: y = 16'hfe01;
			16'he25a: y = 16'hfe01;
			16'he25b: y = 16'hfe01;
			16'he25c: y = 16'hfe01;
			16'he25d: y = 16'hfe01;
			16'he25e: y = 16'hfe01;
			16'he25f: y = 16'hfe01;
			16'he260: y = 16'hfe01;
			16'he261: y = 16'hfe01;
			16'he262: y = 16'hfe01;
			16'he263: y = 16'hfe01;
			16'he264: y = 16'hfe01;
			16'he265: y = 16'hfe01;
			16'he266: y = 16'hfe01;
			16'he267: y = 16'hfe01;
			16'he268: y = 16'hfe01;
			16'he269: y = 16'hfe01;
			16'he26a: y = 16'hfe01;
			16'he26b: y = 16'hfe01;
			16'he26c: y = 16'hfe01;
			16'he26d: y = 16'hfe01;
			16'he26e: y = 16'hfe01;
			16'he26f: y = 16'hfe01;
			16'he270: y = 16'hfe01;
			16'he271: y = 16'hfe01;
			16'he272: y = 16'hfe01;
			16'he273: y = 16'hfe01;
			16'he274: y = 16'hfe01;
			16'he275: y = 16'hfe01;
			16'he276: y = 16'hfe01;
			16'he277: y = 16'hfe01;
			16'he278: y = 16'hfe01;
			16'he279: y = 16'hfe01;
			16'he27a: y = 16'hfe01;
			16'he27b: y = 16'hfe01;
			16'he27c: y = 16'hfe01;
			16'he27d: y = 16'hfe01;
			16'he27e: y = 16'hfe01;
			16'he27f: y = 16'hfe01;
			16'he280: y = 16'hfe01;
			16'he281: y = 16'hfe01;
			16'he282: y = 16'hfe01;
			16'he283: y = 16'hfe01;
			16'he284: y = 16'hfe01;
			16'he285: y = 16'hfe01;
			16'he286: y = 16'hfe01;
			16'he287: y = 16'hfe01;
			16'he288: y = 16'hfe01;
			16'he289: y = 16'hfe01;
			16'he28a: y = 16'hfe01;
			16'he28b: y = 16'hfe01;
			16'he28c: y = 16'hfe01;
			16'he28d: y = 16'hfe01;
			16'he28e: y = 16'hfe01;
			16'he28f: y = 16'hfe01;
			16'he290: y = 16'hfe01;
			16'he291: y = 16'hfe01;
			16'he292: y = 16'hfe01;
			16'he293: y = 16'hfe01;
			16'he294: y = 16'hfe01;
			16'he295: y = 16'hfe01;
			16'he296: y = 16'hfe01;
			16'he297: y = 16'hfe01;
			16'he298: y = 16'hfe01;
			16'he299: y = 16'hfe01;
			16'he29a: y = 16'hfe01;
			16'he29b: y = 16'hfe01;
			16'he29c: y = 16'hfe01;
			16'he29d: y = 16'hfe01;
			16'he29e: y = 16'hfe01;
			16'he29f: y = 16'hfe01;
			16'he2a0: y = 16'hfe01;
			16'he2a1: y = 16'hfe01;
			16'he2a2: y = 16'hfe01;
			16'he2a3: y = 16'hfe01;
			16'he2a4: y = 16'hfe01;
			16'he2a5: y = 16'hfe01;
			16'he2a6: y = 16'hfe01;
			16'he2a7: y = 16'hfe01;
			16'he2a8: y = 16'hfe01;
			16'he2a9: y = 16'hfe01;
			16'he2aa: y = 16'hfe01;
			16'he2ab: y = 16'hfe01;
			16'he2ac: y = 16'hfe01;
			16'he2ad: y = 16'hfe01;
			16'he2ae: y = 16'hfe01;
			16'he2af: y = 16'hfe01;
			16'he2b0: y = 16'hfe01;
			16'he2b1: y = 16'hfe01;
			16'he2b2: y = 16'hfe01;
			16'he2b3: y = 16'hfe01;
			16'he2b4: y = 16'hfe01;
			16'he2b5: y = 16'hfe01;
			16'he2b6: y = 16'hfe01;
			16'he2b7: y = 16'hfe01;
			16'he2b8: y = 16'hfe01;
			16'he2b9: y = 16'hfe01;
			16'he2ba: y = 16'hfe01;
			16'he2bb: y = 16'hfe01;
			16'he2bc: y = 16'hfe01;
			16'he2bd: y = 16'hfe01;
			16'he2be: y = 16'hfe01;
			16'he2bf: y = 16'hfe01;
			16'he2c0: y = 16'hfe01;
			16'he2c1: y = 16'hfe01;
			16'he2c2: y = 16'hfe01;
			16'he2c3: y = 16'hfe01;
			16'he2c4: y = 16'hfe01;
			16'he2c5: y = 16'hfe01;
			16'he2c6: y = 16'hfe01;
			16'he2c7: y = 16'hfe01;
			16'he2c8: y = 16'hfe01;
			16'he2c9: y = 16'hfe01;
			16'he2ca: y = 16'hfe01;
			16'he2cb: y = 16'hfe01;
			16'he2cc: y = 16'hfe01;
			16'he2cd: y = 16'hfe01;
			16'he2ce: y = 16'hfe01;
			16'he2cf: y = 16'hfe01;
			16'he2d0: y = 16'hfe01;
			16'he2d1: y = 16'hfe01;
			16'he2d2: y = 16'hfe01;
			16'he2d3: y = 16'hfe01;
			16'he2d4: y = 16'hfe01;
			16'he2d5: y = 16'hfe01;
			16'he2d6: y = 16'hfe01;
			16'he2d7: y = 16'hfe01;
			16'he2d8: y = 16'hfe01;
			16'he2d9: y = 16'hfe01;
			16'he2da: y = 16'hfe01;
			16'he2db: y = 16'hfe01;
			16'he2dc: y = 16'hfe01;
			16'he2dd: y = 16'hfe01;
			16'he2de: y = 16'hfe01;
			16'he2df: y = 16'hfe01;
			16'he2e0: y = 16'hfe01;
			16'he2e1: y = 16'hfe01;
			16'he2e2: y = 16'hfe01;
			16'he2e3: y = 16'hfe01;
			16'he2e4: y = 16'hfe01;
			16'he2e5: y = 16'hfe01;
			16'he2e6: y = 16'hfe01;
			16'he2e7: y = 16'hfe01;
			16'he2e8: y = 16'hfe01;
			16'he2e9: y = 16'hfe01;
			16'he2ea: y = 16'hfe01;
			16'he2eb: y = 16'hfe01;
			16'he2ec: y = 16'hfe01;
			16'he2ed: y = 16'hfe01;
			16'he2ee: y = 16'hfe01;
			16'he2ef: y = 16'hfe01;
			16'he2f0: y = 16'hfe01;
			16'he2f1: y = 16'hfe01;
			16'he2f2: y = 16'hfe01;
			16'he2f3: y = 16'hfe01;
			16'he2f4: y = 16'hfe01;
			16'he2f5: y = 16'hfe01;
			16'he2f6: y = 16'hfe01;
			16'he2f7: y = 16'hfe01;
			16'he2f8: y = 16'hfe01;
			16'he2f9: y = 16'hfe01;
			16'he2fa: y = 16'hfe01;
			16'he2fb: y = 16'hfe01;
			16'he2fc: y = 16'hfe01;
			16'he2fd: y = 16'hfe01;
			16'he2fe: y = 16'hfe01;
			16'he2ff: y = 16'hfe01;
			16'he300: y = 16'hfe01;
			16'he301: y = 16'hfe01;
			16'he302: y = 16'hfe01;
			16'he303: y = 16'hfe01;
			16'he304: y = 16'hfe01;
			16'he305: y = 16'hfe01;
			16'he306: y = 16'hfe01;
			16'he307: y = 16'hfe01;
			16'he308: y = 16'hfe01;
			16'he309: y = 16'hfe01;
			16'he30a: y = 16'hfe01;
			16'he30b: y = 16'hfe01;
			16'he30c: y = 16'hfe01;
			16'he30d: y = 16'hfe01;
			16'he30e: y = 16'hfe01;
			16'he30f: y = 16'hfe01;
			16'he310: y = 16'hfe01;
			16'he311: y = 16'hfe01;
			16'he312: y = 16'hfe01;
			16'he313: y = 16'hfe01;
			16'he314: y = 16'hfe01;
			16'he315: y = 16'hfe01;
			16'he316: y = 16'hfe01;
			16'he317: y = 16'hfe01;
			16'he318: y = 16'hfe01;
			16'he319: y = 16'hfe01;
			16'he31a: y = 16'hfe01;
			16'he31b: y = 16'hfe01;
			16'he31c: y = 16'hfe01;
			16'he31d: y = 16'hfe01;
			16'he31e: y = 16'hfe01;
			16'he31f: y = 16'hfe01;
			16'he320: y = 16'hfe01;
			16'he321: y = 16'hfe01;
			16'he322: y = 16'hfe01;
			16'he323: y = 16'hfe01;
			16'he324: y = 16'hfe01;
			16'he325: y = 16'hfe01;
			16'he326: y = 16'hfe01;
			16'he327: y = 16'hfe01;
			16'he328: y = 16'hfe01;
			16'he329: y = 16'hfe01;
			16'he32a: y = 16'hfe01;
			16'he32b: y = 16'hfe01;
			16'he32c: y = 16'hfe01;
			16'he32d: y = 16'hfe01;
			16'he32e: y = 16'hfe01;
			16'he32f: y = 16'hfe01;
			16'he330: y = 16'hfe01;
			16'he331: y = 16'hfe01;
			16'he332: y = 16'hfe01;
			16'he333: y = 16'hfe01;
			16'he334: y = 16'hfe01;
			16'he335: y = 16'hfe01;
			16'he336: y = 16'hfe01;
			16'he337: y = 16'hfe01;
			16'he338: y = 16'hfe01;
			16'he339: y = 16'hfe01;
			16'he33a: y = 16'hfe01;
			16'he33b: y = 16'hfe01;
			16'he33c: y = 16'hfe01;
			16'he33d: y = 16'hfe01;
			16'he33e: y = 16'hfe01;
			16'he33f: y = 16'hfe01;
			16'he340: y = 16'hfe01;
			16'he341: y = 16'hfe01;
			16'he342: y = 16'hfe01;
			16'he343: y = 16'hfe01;
			16'he344: y = 16'hfe01;
			16'he345: y = 16'hfe01;
			16'he346: y = 16'hfe01;
			16'he347: y = 16'hfe01;
			16'he348: y = 16'hfe01;
			16'he349: y = 16'hfe01;
			16'he34a: y = 16'hfe01;
			16'he34b: y = 16'hfe01;
			16'he34c: y = 16'hfe01;
			16'he34d: y = 16'hfe01;
			16'he34e: y = 16'hfe01;
			16'he34f: y = 16'hfe01;
			16'he350: y = 16'hfe01;
			16'he351: y = 16'hfe01;
			16'he352: y = 16'hfe01;
			16'he353: y = 16'hfe01;
			16'he354: y = 16'hfe01;
			16'he355: y = 16'hfe01;
			16'he356: y = 16'hfe01;
			16'he357: y = 16'hfe01;
			16'he358: y = 16'hfe01;
			16'he359: y = 16'hfe01;
			16'he35a: y = 16'hfe01;
			16'he35b: y = 16'hfe01;
			16'he35c: y = 16'hfe01;
			16'he35d: y = 16'hfe01;
			16'he35e: y = 16'hfe01;
			16'he35f: y = 16'hfe01;
			16'he360: y = 16'hfe01;
			16'he361: y = 16'hfe01;
			16'he362: y = 16'hfe01;
			16'he363: y = 16'hfe01;
			16'he364: y = 16'hfe01;
			16'he365: y = 16'hfe01;
			16'he366: y = 16'hfe01;
			16'he367: y = 16'hfe01;
			16'he368: y = 16'hfe01;
			16'he369: y = 16'hfe01;
			16'he36a: y = 16'hfe01;
			16'he36b: y = 16'hfe01;
			16'he36c: y = 16'hfe01;
			16'he36d: y = 16'hfe01;
			16'he36e: y = 16'hfe01;
			16'he36f: y = 16'hfe01;
			16'he370: y = 16'hfe01;
			16'he371: y = 16'hfe01;
			16'he372: y = 16'hfe01;
			16'he373: y = 16'hfe01;
			16'he374: y = 16'hfe01;
			16'he375: y = 16'hfe01;
			16'he376: y = 16'hfe01;
			16'he377: y = 16'hfe01;
			16'he378: y = 16'hfe01;
			16'he379: y = 16'hfe01;
			16'he37a: y = 16'hfe01;
			16'he37b: y = 16'hfe01;
			16'he37c: y = 16'hfe01;
			16'he37d: y = 16'hfe01;
			16'he37e: y = 16'hfe01;
			16'he37f: y = 16'hfe01;
			16'he380: y = 16'hfe01;
			16'he381: y = 16'hfe01;
			16'he382: y = 16'hfe01;
			16'he383: y = 16'hfe01;
			16'he384: y = 16'hfe01;
			16'he385: y = 16'hfe01;
			16'he386: y = 16'hfe01;
			16'he387: y = 16'hfe01;
			16'he388: y = 16'hfe01;
			16'he389: y = 16'hfe01;
			16'he38a: y = 16'hfe01;
			16'he38b: y = 16'hfe01;
			16'he38c: y = 16'hfe01;
			16'he38d: y = 16'hfe01;
			16'he38e: y = 16'hfe01;
			16'he38f: y = 16'hfe01;
			16'he390: y = 16'hfe01;
			16'he391: y = 16'hfe01;
			16'he392: y = 16'hfe01;
			16'he393: y = 16'hfe01;
			16'he394: y = 16'hfe01;
			16'he395: y = 16'hfe01;
			16'he396: y = 16'hfe01;
			16'he397: y = 16'hfe01;
			16'he398: y = 16'hfe01;
			16'he399: y = 16'hfe01;
			16'he39a: y = 16'hfe01;
			16'he39b: y = 16'hfe01;
			16'he39c: y = 16'hfe01;
			16'he39d: y = 16'hfe01;
			16'he39e: y = 16'hfe01;
			16'he39f: y = 16'hfe01;
			16'he3a0: y = 16'hfe01;
			16'he3a1: y = 16'hfe01;
			16'he3a2: y = 16'hfe01;
			16'he3a3: y = 16'hfe01;
			16'he3a4: y = 16'hfe01;
			16'he3a5: y = 16'hfe01;
			16'he3a6: y = 16'hfe01;
			16'he3a7: y = 16'hfe01;
			16'he3a8: y = 16'hfe01;
			16'he3a9: y = 16'hfe01;
			16'he3aa: y = 16'hfe01;
			16'he3ab: y = 16'hfe01;
			16'he3ac: y = 16'hfe01;
			16'he3ad: y = 16'hfe01;
			16'he3ae: y = 16'hfe01;
			16'he3af: y = 16'hfe01;
			16'he3b0: y = 16'hfe01;
			16'he3b1: y = 16'hfe01;
			16'he3b2: y = 16'hfe01;
			16'he3b3: y = 16'hfe01;
			16'he3b4: y = 16'hfe01;
			16'he3b5: y = 16'hfe01;
			16'he3b6: y = 16'hfe01;
			16'he3b7: y = 16'hfe01;
			16'he3b8: y = 16'hfe01;
			16'he3b9: y = 16'hfe01;
			16'he3ba: y = 16'hfe01;
			16'he3bb: y = 16'hfe01;
			16'he3bc: y = 16'hfe01;
			16'he3bd: y = 16'hfe01;
			16'he3be: y = 16'hfe01;
			16'he3bf: y = 16'hfe01;
			16'he3c0: y = 16'hfe01;
			16'he3c1: y = 16'hfe01;
			16'he3c2: y = 16'hfe01;
			16'he3c3: y = 16'hfe01;
			16'he3c4: y = 16'hfe01;
			16'he3c5: y = 16'hfe01;
			16'he3c6: y = 16'hfe01;
			16'he3c7: y = 16'hfe01;
			16'he3c8: y = 16'hfe01;
			16'he3c9: y = 16'hfe01;
			16'he3ca: y = 16'hfe01;
			16'he3cb: y = 16'hfe01;
			16'he3cc: y = 16'hfe01;
			16'he3cd: y = 16'hfe01;
			16'he3ce: y = 16'hfe01;
			16'he3cf: y = 16'hfe01;
			16'he3d0: y = 16'hfe01;
			16'he3d1: y = 16'hfe01;
			16'he3d2: y = 16'hfe01;
			16'he3d3: y = 16'hfe01;
			16'he3d4: y = 16'hfe01;
			16'he3d5: y = 16'hfe01;
			16'he3d6: y = 16'hfe01;
			16'he3d7: y = 16'hfe01;
			16'he3d8: y = 16'hfe01;
			16'he3d9: y = 16'hfe01;
			16'he3da: y = 16'hfe01;
			16'he3db: y = 16'hfe01;
			16'he3dc: y = 16'hfe01;
			16'he3dd: y = 16'hfe01;
			16'he3de: y = 16'hfe01;
			16'he3df: y = 16'hfe01;
			16'he3e0: y = 16'hfe01;
			16'he3e1: y = 16'hfe01;
			16'he3e2: y = 16'hfe01;
			16'he3e3: y = 16'hfe01;
			16'he3e4: y = 16'hfe01;
			16'he3e5: y = 16'hfe01;
			16'he3e6: y = 16'hfe01;
			16'he3e7: y = 16'hfe01;
			16'he3e8: y = 16'hfe01;
			16'he3e9: y = 16'hfe01;
			16'he3ea: y = 16'hfe01;
			16'he3eb: y = 16'hfe01;
			16'he3ec: y = 16'hfe01;
			16'he3ed: y = 16'hfe01;
			16'he3ee: y = 16'hfe01;
			16'he3ef: y = 16'hfe01;
			16'he3f0: y = 16'hfe01;
			16'he3f1: y = 16'hfe01;
			16'he3f2: y = 16'hfe01;
			16'he3f3: y = 16'hfe01;
			16'he3f4: y = 16'hfe01;
			16'he3f5: y = 16'hfe01;
			16'he3f6: y = 16'hfe01;
			16'he3f7: y = 16'hfe01;
			16'he3f8: y = 16'hfe01;
			16'he3f9: y = 16'hfe01;
			16'he3fa: y = 16'hfe01;
			16'he3fb: y = 16'hfe01;
			16'he3fc: y = 16'hfe01;
			16'he3fd: y = 16'hfe01;
			16'he3fe: y = 16'hfe01;
			16'he3ff: y = 16'hfe01;
			16'he400: y = 16'hfe01;
			16'he401: y = 16'hfe01;
			16'he402: y = 16'hfe01;
			16'he403: y = 16'hfe01;
			16'he404: y = 16'hfe01;
			16'he405: y = 16'hfe01;
			16'he406: y = 16'hfe01;
			16'he407: y = 16'hfe01;
			16'he408: y = 16'hfe01;
			16'he409: y = 16'hfe01;
			16'he40a: y = 16'hfe01;
			16'he40b: y = 16'hfe01;
			16'he40c: y = 16'hfe01;
			16'he40d: y = 16'hfe01;
			16'he40e: y = 16'hfe01;
			16'he40f: y = 16'hfe01;
			16'he410: y = 16'hfe01;
			16'he411: y = 16'hfe01;
			16'he412: y = 16'hfe01;
			16'he413: y = 16'hfe01;
			16'he414: y = 16'hfe01;
			16'he415: y = 16'hfe01;
			16'he416: y = 16'hfe01;
			16'he417: y = 16'hfe01;
			16'he418: y = 16'hfe01;
			16'he419: y = 16'hfe01;
			16'he41a: y = 16'hfe01;
			16'he41b: y = 16'hfe01;
			16'he41c: y = 16'hfe01;
			16'he41d: y = 16'hfe01;
			16'he41e: y = 16'hfe01;
			16'he41f: y = 16'hfe01;
			16'he420: y = 16'hfe01;
			16'he421: y = 16'hfe01;
			16'he422: y = 16'hfe01;
			16'he423: y = 16'hfe01;
			16'he424: y = 16'hfe01;
			16'he425: y = 16'hfe01;
			16'he426: y = 16'hfe01;
			16'he427: y = 16'hfe01;
			16'he428: y = 16'hfe01;
			16'he429: y = 16'hfe01;
			16'he42a: y = 16'hfe01;
			16'he42b: y = 16'hfe01;
			16'he42c: y = 16'hfe01;
			16'he42d: y = 16'hfe01;
			16'he42e: y = 16'hfe01;
			16'he42f: y = 16'hfe01;
			16'he430: y = 16'hfe01;
			16'he431: y = 16'hfe01;
			16'he432: y = 16'hfe01;
			16'he433: y = 16'hfe01;
			16'he434: y = 16'hfe01;
			16'he435: y = 16'hfe01;
			16'he436: y = 16'hfe01;
			16'he437: y = 16'hfe01;
			16'he438: y = 16'hfe01;
			16'he439: y = 16'hfe01;
			16'he43a: y = 16'hfe01;
			16'he43b: y = 16'hfe01;
			16'he43c: y = 16'hfe01;
			16'he43d: y = 16'hfe01;
			16'he43e: y = 16'hfe01;
			16'he43f: y = 16'hfe01;
			16'he440: y = 16'hfe01;
			16'he441: y = 16'hfe01;
			16'he442: y = 16'hfe01;
			16'he443: y = 16'hfe01;
			16'he444: y = 16'hfe01;
			16'he445: y = 16'hfe01;
			16'he446: y = 16'hfe01;
			16'he447: y = 16'hfe01;
			16'he448: y = 16'hfe01;
			16'he449: y = 16'hfe01;
			16'he44a: y = 16'hfe01;
			16'he44b: y = 16'hfe01;
			16'he44c: y = 16'hfe01;
			16'he44d: y = 16'hfe01;
			16'he44e: y = 16'hfe01;
			16'he44f: y = 16'hfe01;
			16'he450: y = 16'hfe01;
			16'he451: y = 16'hfe01;
			16'he452: y = 16'hfe01;
			16'he453: y = 16'hfe01;
			16'he454: y = 16'hfe01;
			16'he455: y = 16'hfe01;
			16'he456: y = 16'hfe01;
			16'he457: y = 16'hfe01;
			16'he458: y = 16'hfe01;
			16'he459: y = 16'hfe01;
			16'he45a: y = 16'hfe01;
			16'he45b: y = 16'hfe01;
			16'he45c: y = 16'hfe01;
			16'he45d: y = 16'hfe01;
			16'he45e: y = 16'hfe01;
			16'he45f: y = 16'hfe01;
			16'he460: y = 16'hfe01;
			16'he461: y = 16'hfe01;
			16'he462: y = 16'hfe01;
			16'he463: y = 16'hfe01;
			16'he464: y = 16'hfe01;
			16'he465: y = 16'hfe01;
			16'he466: y = 16'hfe01;
			16'he467: y = 16'hfe01;
			16'he468: y = 16'hfe01;
			16'he469: y = 16'hfe01;
			16'he46a: y = 16'hfe01;
			16'he46b: y = 16'hfe01;
			16'he46c: y = 16'hfe01;
			16'he46d: y = 16'hfe01;
			16'he46e: y = 16'hfe01;
			16'he46f: y = 16'hfe01;
			16'he470: y = 16'hfe01;
			16'he471: y = 16'hfe01;
			16'he472: y = 16'hfe01;
			16'he473: y = 16'hfe01;
			16'he474: y = 16'hfe01;
			16'he475: y = 16'hfe01;
			16'he476: y = 16'hfe01;
			16'he477: y = 16'hfe01;
			16'he478: y = 16'hfe01;
			16'he479: y = 16'hfe01;
			16'he47a: y = 16'hfe01;
			16'he47b: y = 16'hfe01;
			16'he47c: y = 16'hfe01;
			16'he47d: y = 16'hfe01;
			16'he47e: y = 16'hfe01;
			16'he47f: y = 16'hfe01;
			16'he480: y = 16'hfe01;
			16'he481: y = 16'hfe01;
			16'he482: y = 16'hfe01;
			16'he483: y = 16'hfe01;
			16'he484: y = 16'hfe01;
			16'he485: y = 16'hfe01;
			16'he486: y = 16'hfe01;
			16'he487: y = 16'hfe01;
			16'he488: y = 16'hfe01;
			16'he489: y = 16'hfe01;
			16'he48a: y = 16'hfe01;
			16'he48b: y = 16'hfe01;
			16'he48c: y = 16'hfe01;
			16'he48d: y = 16'hfe01;
			16'he48e: y = 16'hfe01;
			16'he48f: y = 16'hfe01;
			16'he490: y = 16'hfe01;
			16'he491: y = 16'hfe01;
			16'he492: y = 16'hfe01;
			16'he493: y = 16'hfe01;
			16'he494: y = 16'hfe01;
			16'he495: y = 16'hfe01;
			16'he496: y = 16'hfe01;
			16'he497: y = 16'hfe01;
			16'he498: y = 16'hfe01;
			16'he499: y = 16'hfe01;
			16'he49a: y = 16'hfe01;
			16'he49b: y = 16'hfe01;
			16'he49c: y = 16'hfe01;
			16'he49d: y = 16'hfe01;
			16'he49e: y = 16'hfe01;
			16'he49f: y = 16'hfe01;
			16'he4a0: y = 16'hfe01;
			16'he4a1: y = 16'hfe01;
			16'he4a2: y = 16'hfe01;
			16'he4a3: y = 16'hfe01;
			16'he4a4: y = 16'hfe01;
			16'he4a5: y = 16'hfe01;
			16'he4a6: y = 16'hfe01;
			16'he4a7: y = 16'hfe01;
			16'he4a8: y = 16'hfe01;
			16'he4a9: y = 16'hfe01;
			16'he4aa: y = 16'hfe01;
			16'he4ab: y = 16'hfe01;
			16'he4ac: y = 16'hfe01;
			16'he4ad: y = 16'hfe01;
			16'he4ae: y = 16'hfe01;
			16'he4af: y = 16'hfe01;
			16'he4b0: y = 16'hfe01;
			16'he4b1: y = 16'hfe01;
			16'he4b2: y = 16'hfe01;
			16'he4b3: y = 16'hfe01;
			16'he4b4: y = 16'hfe01;
			16'he4b5: y = 16'hfe01;
			16'he4b6: y = 16'hfe01;
			16'he4b7: y = 16'hfe01;
			16'he4b8: y = 16'hfe01;
			16'he4b9: y = 16'hfe01;
			16'he4ba: y = 16'hfe01;
			16'he4bb: y = 16'hfe01;
			16'he4bc: y = 16'hfe01;
			16'he4bd: y = 16'hfe01;
			16'he4be: y = 16'hfe01;
			16'he4bf: y = 16'hfe01;
			16'he4c0: y = 16'hfe01;
			16'he4c1: y = 16'hfe01;
			16'he4c2: y = 16'hfe01;
			16'he4c3: y = 16'hfe01;
			16'he4c4: y = 16'hfe01;
			16'he4c5: y = 16'hfe01;
			16'he4c6: y = 16'hfe01;
			16'he4c7: y = 16'hfe01;
			16'he4c8: y = 16'hfe01;
			16'he4c9: y = 16'hfe01;
			16'he4ca: y = 16'hfe01;
			16'he4cb: y = 16'hfe01;
			16'he4cc: y = 16'hfe01;
			16'he4cd: y = 16'hfe01;
			16'he4ce: y = 16'hfe01;
			16'he4cf: y = 16'hfe01;
			16'he4d0: y = 16'hfe01;
			16'he4d1: y = 16'hfe01;
			16'he4d2: y = 16'hfe01;
			16'he4d3: y = 16'hfe01;
			16'he4d4: y = 16'hfe01;
			16'he4d5: y = 16'hfe01;
			16'he4d6: y = 16'hfe01;
			16'he4d7: y = 16'hfe01;
			16'he4d8: y = 16'hfe01;
			16'he4d9: y = 16'hfe01;
			16'he4da: y = 16'hfe01;
			16'he4db: y = 16'hfe01;
			16'he4dc: y = 16'hfe01;
			16'he4dd: y = 16'hfe01;
			16'he4de: y = 16'hfe01;
			16'he4df: y = 16'hfe01;
			16'he4e0: y = 16'hfe01;
			16'he4e1: y = 16'hfe01;
			16'he4e2: y = 16'hfe01;
			16'he4e3: y = 16'hfe01;
			16'he4e4: y = 16'hfe01;
			16'he4e5: y = 16'hfe01;
			16'he4e6: y = 16'hfe01;
			16'he4e7: y = 16'hfe01;
			16'he4e8: y = 16'hfe01;
			16'he4e9: y = 16'hfe01;
			16'he4ea: y = 16'hfe01;
			16'he4eb: y = 16'hfe01;
			16'he4ec: y = 16'hfe01;
			16'he4ed: y = 16'hfe01;
			16'he4ee: y = 16'hfe01;
			16'he4ef: y = 16'hfe01;
			16'he4f0: y = 16'hfe01;
			16'he4f1: y = 16'hfe01;
			16'he4f2: y = 16'hfe01;
			16'he4f3: y = 16'hfe01;
			16'he4f4: y = 16'hfe01;
			16'he4f5: y = 16'hfe01;
			16'he4f6: y = 16'hfe01;
			16'he4f7: y = 16'hfe01;
			16'he4f8: y = 16'hfe01;
			16'he4f9: y = 16'hfe01;
			16'he4fa: y = 16'hfe01;
			16'he4fb: y = 16'hfe01;
			16'he4fc: y = 16'hfe01;
			16'he4fd: y = 16'hfe01;
			16'he4fe: y = 16'hfe01;
			16'he4ff: y = 16'hfe01;
			16'he500: y = 16'hfe01;
			16'he501: y = 16'hfe01;
			16'he502: y = 16'hfe01;
			16'he503: y = 16'hfe01;
			16'he504: y = 16'hfe01;
			16'he505: y = 16'hfe01;
			16'he506: y = 16'hfe01;
			16'he507: y = 16'hfe01;
			16'he508: y = 16'hfe01;
			16'he509: y = 16'hfe01;
			16'he50a: y = 16'hfe01;
			16'he50b: y = 16'hfe01;
			16'he50c: y = 16'hfe01;
			16'he50d: y = 16'hfe01;
			16'he50e: y = 16'hfe01;
			16'he50f: y = 16'hfe01;
			16'he510: y = 16'hfe01;
			16'he511: y = 16'hfe01;
			16'he512: y = 16'hfe01;
			16'he513: y = 16'hfe01;
			16'he514: y = 16'hfe01;
			16'he515: y = 16'hfe01;
			16'he516: y = 16'hfe01;
			16'he517: y = 16'hfe01;
			16'he518: y = 16'hfe01;
			16'he519: y = 16'hfe01;
			16'he51a: y = 16'hfe01;
			16'he51b: y = 16'hfe01;
			16'he51c: y = 16'hfe01;
			16'he51d: y = 16'hfe01;
			16'he51e: y = 16'hfe01;
			16'he51f: y = 16'hfe01;
			16'he520: y = 16'hfe01;
			16'he521: y = 16'hfe01;
			16'he522: y = 16'hfe01;
			16'he523: y = 16'hfe01;
			16'he524: y = 16'hfe01;
			16'he525: y = 16'hfe01;
			16'he526: y = 16'hfe01;
			16'he527: y = 16'hfe01;
			16'he528: y = 16'hfe01;
			16'he529: y = 16'hfe01;
			16'he52a: y = 16'hfe01;
			16'he52b: y = 16'hfe01;
			16'he52c: y = 16'hfe01;
			16'he52d: y = 16'hfe01;
			16'he52e: y = 16'hfe01;
			16'he52f: y = 16'hfe01;
			16'he530: y = 16'hfe01;
			16'he531: y = 16'hfe01;
			16'he532: y = 16'hfe01;
			16'he533: y = 16'hfe01;
			16'he534: y = 16'hfe01;
			16'he535: y = 16'hfe01;
			16'he536: y = 16'hfe01;
			16'he537: y = 16'hfe01;
			16'he538: y = 16'hfe01;
			16'he539: y = 16'hfe01;
			16'he53a: y = 16'hfe01;
			16'he53b: y = 16'hfe01;
			16'he53c: y = 16'hfe01;
			16'he53d: y = 16'hfe01;
			16'he53e: y = 16'hfe01;
			16'he53f: y = 16'hfe01;
			16'he540: y = 16'hfe01;
			16'he541: y = 16'hfe01;
			16'he542: y = 16'hfe01;
			16'he543: y = 16'hfe01;
			16'he544: y = 16'hfe01;
			16'he545: y = 16'hfe01;
			16'he546: y = 16'hfe01;
			16'he547: y = 16'hfe01;
			16'he548: y = 16'hfe01;
			16'he549: y = 16'hfe01;
			16'he54a: y = 16'hfe01;
			16'he54b: y = 16'hfe01;
			16'he54c: y = 16'hfe01;
			16'he54d: y = 16'hfe01;
			16'he54e: y = 16'hfe01;
			16'he54f: y = 16'hfe01;
			16'he550: y = 16'hfe01;
			16'he551: y = 16'hfe01;
			16'he552: y = 16'hfe01;
			16'he553: y = 16'hfe01;
			16'he554: y = 16'hfe01;
			16'he555: y = 16'hfe01;
			16'he556: y = 16'hfe01;
			16'he557: y = 16'hfe01;
			16'he558: y = 16'hfe01;
			16'he559: y = 16'hfe01;
			16'he55a: y = 16'hfe01;
			16'he55b: y = 16'hfe01;
			16'he55c: y = 16'hfe01;
			16'he55d: y = 16'hfe01;
			16'he55e: y = 16'hfe01;
			16'he55f: y = 16'hfe01;
			16'he560: y = 16'hfe01;
			16'he561: y = 16'hfe01;
			16'he562: y = 16'hfe01;
			16'he563: y = 16'hfe01;
			16'he564: y = 16'hfe01;
			16'he565: y = 16'hfe01;
			16'he566: y = 16'hfe01;
			16'he567: y = 16'hfe01;
			16'he568: y = 16'hfe01;
			16'he569: y = 16'hfe01;
			16'he56a: y = 16'hfe01;
			16'he56b: y = 16'hfe01;
			16'he56c: y = 16'hfe01;
			16'he56d: y = 16'hfe01;
			16'he56e: y = 16'hfe01;
			16'he56f: y = 16'hfe01;
			16'he570: y = 16'hfe01;
			16'he571: y = 16'hfe01;
			16'he572: y = 16'hfe01;
			16'he573: y = 16'hfe01;
			16'he574: y = 16'hfe01;
			16'he575: y = 16'hfe01;
			16'he576: y = 16'hfe01;
			16'he577: y = 16'hfe01;
			16'he578: y = 16'hfe01;
			16'he579: y = 16'hfe01;
			16'he57a: y = 16'hfe01;
			16'he57b: y = 16'hfe01;
			16'he57c: y = 16'hfe01;
			16'he57d: y = 16'hfe01;
			16'he57e: y = 16'hfe01;
			16'he57f: y = 16'hfe01;
			16'he580: y = 16'hfe01;
			16'he581: y = 16'hfe01;
			16'he582: y = 16'hfe01;
			16'he583: y = 16'hfe01;
			16'he584: y = 16'hfe01;
			16'he585: y = 16'hfe01;
			16'he586: y = 16'hfe01;
			16'he587: y = 16'hfe01;
			16'he588: y = 16'hfe01;
			16'he589: y = 16'hfe01;
			16'he58a: y = 16'hfe01;
			16'he58b: y = 16'hfe01;
			16'he58c: y = 16'hfe01;
			16'he58d: y = 16'hfe01;
			16'he58e: y = 16'hfe01;
			16'he58f: y = 16'hfe01;
			16'he590: y = 16'hfe01;
			16'he591: y = 16'hfe01;
			16'he592: y = 16'hfe01;
			16'he593: y = 16'hfe01;
			16'he594: y = 16'hfe01;
			16'he595: y = 16'hfe01;
			16'he596: y = 16'hfe01;
			16'he597: y = 16'hfe01;
			16'he598: y = 16'hfe01;
			16'he599: y = 16'hfe01;
			16'he59a: y = 16'hfe01;
			16'he59b: y = 16'hfe01;
			16'he59c: y = 16'hfe01;
			16'he59d: y = 16'hfe01;
			16'he59e: y = 16'hfe01;
			16'he59f: y = 16'hfe01;
			16'he5a0: y = 16'hfe01;
			16'he5a1: y = 16'hfe01;
			16'he5a2: y = 16'hfe01;
			16'he5a3: y = 16'hfe01;
			16'he5a4: y = 16'hfe01;
			16'he5a5: y = 16'hfe01;
			16'he5a6: y = 16'hfe01;
			16'he5a7: y = 16'hfe01;
			16'he5a8: y = 16'hfe01;
			16'he5a9: y = 16'hfe01;
			16'he5aa: y = 16'hfe01;
			16'he5ab: y = 16'hfe01;
			16'he5ac: y = 16'hfe01;
			16'he5ad: y = 16'hfe01;
			16'he5ae: y = 16'hfe01;
			16'he5af: y = 16'hfe01;
			16'he5b0: y = 16'hfe01;
			16'he5b1: y = 16'hfe01;
			16'he5b2: y = 16'hfe01;
			16'he5b3: y = 16'hfe01;
			16'he5b4: y = 16'hfe01;
			16'he5b5: y = 16'hfe01;
			16'he5b6: y = 16'hfe01;
			16'he5b7: y = 16'hfe01;
			16'he5b8: y = 16'hfe01;
			16'he5b9: y = 16'hfe01;
			16'he5ba: y = 16'hfe01;
			16'he5bb: y = 16'hfe01;
			16'he5bc: y = 16'hfe01;
			16'he5bd: y = 16'hfe01;
			16'he5be: y = 16'hfe01;
			16'he5bf: y = 16'hfe01;
			16'he5c0: y = 16'hfe01;
			16'he5c1: y = 16'hfe01;
			16'he5c2: y = 16'hfe01;
			16'he5c3: y = 16'hfe01;
			16'he5c4: y = 16'hfe01;
			16'he5c5: y = 16'hfe01;
			16'he5c6: y = 16'hfe01;
			16'he5c7: y = 16'hfe01;
			16'he5c8: y = 16'hfe01;
			16'he5c9: y = 16'hfe01;
			16'he5ca: y = 16'hfe01;
			16'he5cb: y = 16'hfe01;
			16'he5cc: y = 16'hfe01;
			16'he5cd: y = 16'hfe01;
			16'he5ce: y = 16'hfe01;
			16'he5cf: y = 16'hfe01;
			16'he5d0: y = 16'hfe01;
			16'he5d1: y = 16'hfe01;
			16'he5d2: y = 16'hfe01;
			16'he5d3: y = 16'hfe01;
			16'he5d4: y = 16'hfe01;
			16'he5d5: y = 16'hfe01;
			16'he5d6: y = 16'hfe01;
			16'he5d7: y = 16'hfe01;
			16'he5d8: y = 16'hfe01;
			16'he5d9: y = 16'hfe01;
			16'he5da: y = 16'hfe01;
			16'he5db: y = 16'hfe01;
			16'he5dc: y = 16'hfe01;
			16'he5dd: y = 16'hfe01;
			16'he5de: y = 16'hfe01;
			16'he5df: y = 16'hfe01;
			16'he5e0: y = 16'hfe01;
			16'he5e1: y = 16'hfe01;
			16'he5e2: y = 16'hfe01;
			16'he5e3: y = 16'hfe01;
			16'he5e4: y = 16'hfe01;
			16'he5e5: y = 16'hfe01;
			16'he5e6: y = 16'hfe01;
			16'he5e7: y = 16'hfe01;
			16'he5e8: y = 16'hfe01;
			16'he5e9: y = 16'hfe01;
			16'he5ea: y = 16'hfe01;
			16'he5eb: y = 16'hfe01;
			16'he5ec: y = 16'hfe01;
			16'he5ed: y = 16'hfe01;
			16'he5ee: y = 16'hfe01;
			16'he5ef: y = 16'hfe01;
			16'he5f0: y = 16'hfe01;
			16'he5f1: y = 16'hfe01;
			16'he5f2: y = 16'hfe01;
			16'he5f3: y = 16'hfe01;
			16'he5f4: y = 16'hfe01;
			16'he5f5: y = 16'hfe01;
			16'he5f6: y = 16'hfe01;
			16'he5f7: y = 16'hfe01;
			16'he5f8: y = 16'hfe01;
			16'he5f9: y = 16'hfe01;
			16'he5fa: y = 16'hfe01;
			16'he5fb: y = 16'hfe01;
			16'he5fc: y = 16'hfe01;
			16'he5fd: y = 16'hfe01;
			16'he5fe: y = 16'hfe01;
			16'he5ff: y = 16'hfe01;
			16'he600: y = 16'hfe01;
			16'he601: y = 16'hfe01;
			16'he602: y = 16'hfe01;
			16'he603: y = 16'hfe01;
			16'he604: y = 16'hfe01;
			16'he605: y = 16'hfe01;
			16'he606: y = 16'hfe01;
			16'he607: y = 16'hfe01;
			16'he608: y = 16'hfe01;
			16'he609: y = 16'hfe01;
			16'he60a: y = 16'hfe01;
			16'he60b: y = 16'hfe01;
			16'he60c: y = 16'hfe01;
			16'he60d: y = 16'hfe01;
			16'he60e: y = 16'hfe01;
			16'he60f: y = 16'hfe01;
			16'he610: y = 16'hfe01;
			16'he611: y = 16'hfe01;
			16'he612: y = 16'hfe01;
			16'he613: y = 16'hfe01;
			16'he614: y = 16'hfe01;
			16'he615: y = 16'hfe01;
			16'he616: y = 16'hfe01;
			16'he617: y = 16'hfe01;
			16'he618: y = 16'hfe01;
			16'he619: y = 16'hfe01;
			16'he61a: y = 16'hfe01;
			16'he61b: y = 16'hfe01;
			16'he61c: y = 16'hfe01;
			16'he61d: y = 16'hfe01;
			16'he61e: y = 16'hfe01;
			16'he61f: y = 16'hfe01;
			16'he620: y = 16'hfe01;
			16'he621: y = 16'hfe01;
			16'he622: y = 16'hfe01;
			16'he623: y = 16'hfe01;
			16'he624: y = 16'hfe01;
			16'he625: y = 16'hfe01;
			16'he626: y = 16'hfe01;
			16'he627: y = 16'hfe01;
			16'he628: y = 16'hfe01;
			16'he629: y = 16'hfe01;
			16'he62a: y = 16'hfe01;
			16'he62b: y = 16'hfe01;
			16'he62c: y = 16'hfe01;
			16'he62d: y = 16'hfe01;
			16'he62e: y = 16'hfe01;
			16'he62f: y = 16'hfe01;
			16'he630: y = 16'hfe01;
			16'he631: y = 16'hfe01;
			16'he632: y = 16'hfe01;
			16'he633: y = 16'hfe01;
			16'he634: y = 16'hfe01;
			16'he635: y = 16'hfe01;
			16'he636: y = 16'hfe01;
			16'he637: y = 16'hfe01;
			16'he638: y = 16'hfe01;
			16'he639: y = 16'hfe01;
			16'he63a: y = 16'hfe01;
			16'he63b: y = 16'hfe01;
			16'he63c: y = 16'hfe01;
			16'he63d: y = 16'hfe01;
			16'he63e: y = 16'hfe01;
			16'he63f: y = 16'hfe01;
			16'he640: y = 16'hfe01;
			16'he641: y = 16'hfe01;
			16'he642: y = 16'hfe01;
			16'he643: y = 16'hfe01;
			16'he644: y = 16'hfe01;
			16'he645: y = 16'hfe01;
			16'he646: y = 16'hfe01;
			16'he647: y = 16'hfe01;
			16'he648: y = 16'hfe01;
			16'he649: y = 16'hfe01;
			16'he64a: y = 16'hfe01;
			16'he64b: y = 16'hfe01;
			16'he64c: y = 16'hfe01;
			16'he64d: y = 16'hfe01;
			16'he64e: y = 16'hfe01;
			16'he64f: y = 16'hfe01;
			16'he650: y = 16'hfe01;
			16'he651: y = 16'hfe01;
			16'he652: y = 16'hfe01;
			16'he653: y = 16'hfe01;
			16'he654: y = 16'hfe01;
			16'he655: y = 16'hfe01;
			16'he656: y = 16'hfe01;
			16'he657: y = 16'hfe01;
			16'he658: y = 16'hfe01;
			16'he659: y = 16'hfe01;
			16'he65a: y = 16'hfe01;
			16'he65b: y = 16'hfe01;
			16'he65c: y = 16'hfe01;
			16'he65d: y = 16'hfe01;
			16'he65e: y = 16'hfe01;
			16'he65f: y = 16'hfe01;
			16'he660: y = 16'hfe01;
			16'he661: y = 16'hfe01;
			16'he662: y = 16'hfe01;
			16'he663: y = 16'hfe01;
			16'he664: y = 16'hfe01;
			16'he665: y = 16'hfe01;
			16'he666: y = 16'hfe01;
			16'he667: y = 16'hfe01;
			16'he668: y = 16'hfe01;
			16'he669: y = 16'hfe01;
			16'he66a: y = 16'hfe01;
			16'he66b: y = 16'hfe01;
			16'he66c: y = 16'hfe01;
			16'he66d: y = 16'hfe01;
			16'he66e: y = 16'hfe01;
			16'he66f: y = 16'hfe01;
			16'he670: y = 16'hfe01;
			16'he671: y = 16'hfe01;
			16'he672: y = 16'hfe01;
			16'he673: y = 16'hfe01;
			16'he674: y = 16'hfe01;
			16'he675: y = 16'hfe01;
			16'he676: y = 16'hfe01;
			16'he677: y = 16'hfe01;
			16'he678: y = 16'hfe01;
			16'he679: y = 16'hfe01;
			16'he67a: y = 16'hfe01;
			16'he67b: y = 16'hfe01;
			16'he67c: y = 16'hfe01;
			16'he67d: y = 16'hfe01;
			16'he67e: y = 16'hfe01;
			16'he67f: y = 16'hfe01;
			16'he680: y = 16'hfe01;
			16'he681: y = 16'hfe01;
			16'he682: y = 16'hfe01;
			16'he683: y = 16'hfe01;
			16'he684: y = 16'hfe01;
			16'he685: y = 16'hfe01;
			16'he686: y = 16'hfe01;
			16'he687: y = 16'hfe01;
			16'he688: y = 16'hfe01;
			16'he689: y = 16'hfe01;
			16'he68a: y = 16'hfe01;
			16'he68b: y = 16'hfe01;
			16'he68c: y = 16'hfe01;
			16'he68d: y = 16'hfe01;
			16'he68e: y = 16'hfe01;
			16'he68f: y = 16'hfe01;
			16'he690: y = 16'hfe01;
			16'he691: y = 16'hfe01;
			16'he692: y = 16'hfe01;
			16'he693: y = 16'hfe01;
			16'he694: y = 16'hfe01;
			16'he695: y = 16'hfe01;
			16'he696: y = 16'hfe01;
			16'he697: y = 16'hfe01;
			16'he698: y = 16'hfe01;
			16'he699: y = 16'hfe01;
			16'he69a: y = 16'hfe01;
			16'he69b: y = 16'hfe01;
			16'he69c: y = 16'hfe01;
			16'he69d: y = 16'hfe01;
			16'he69e: y = 16'hfe01;
			16'he69f: y = 16'hfe01;
			16'he6a0: y = 16'hfe01;
			16'he6a1: y = 16'hfe01;
			16'he6a2: y = 16'hfe01;
			16'he6a3: y = 16'hfe01;
			16'he6a4: y = 16'hfe01;
			16'he6a5: y = 16'hfe01;
			16'he6a6: y = 16'hfe01;
			16'he6a7: y = 16'hfe01;
			16'he6a8: y = 16'hfe01;
			16'he6a9: y = 16'hfe01;
			16'he6aa: y = 16'hfe01;
			16'he6ab: y = 16'hfe01;
			16'he6ac: y = 16'hfe01;
			16'he6ad: y = 16'hfe01;
			16'he6ae: y = 16'hfe01;
			16'he6af: y = 16'hfe01;
			16'he6b0: y = 16'hfe01;
			16'he6b1: y = 16'hfe01;
			16'he6b2: y = 16'hfe01;
			16'he6b3: y = 16'hfe01;
			16'he6b4: y = 16'hfe01;
			16'he6b5: y = 16'hfe01;
			16'he6b6: y = 16'hfe01;
			16'he6b7: y = 16'hfe01;
			16'he6b8: y = 16'hfe01;
			16'he6b9: y = 16'hfe01;
			16'he6ba: y = 16'hfe01;
			16'he6bb: y = 16'hfe01;
			16'he6bc: y = 16'hfe01;
			16'he6bd: y = 16'hfe01;
			16'he6be: y = 16'hfe01;
			16'he6bf: y = 16'hfe01;
			16'he6c0: y = 16'hfe01;
			16'he6c1: y = 16'hfe01;
			16'he6c2: y = 16'hfe01;
			16'he6c3: y = 16'hfe01;
			16'he6c4: y = 16'hfe01;
			16'he6c5: y = 16'hfe01;
			16'he6c6: y = 16'hfe01;
			16'he6c7: y = 16'hfe01;
			16'he6c8: y = 16'hfe01;
			16'he6c9: y = 16'hfe01;
			16'he6ca: y = 16'hfe01;
			16'he6cb: y = 16'hfe01;
			16'he6cc: y = 16'hfe01;
			16'he6cd: y = 16'hfe01;
			16'he6ce: y = 16'hfe01;
			16'he6cf: y = 16'hfe01;
			16'he6d0: y = 16'hfe01;
			16'he6d1: y = 16'hfe01;
			16'he6d2: y = 16'hfe01;
			16'he6d3: y = 16'hfe01;
			16'he6d4: y = 16'hfe01;
			16'he6d5: y = 16'hfe01;
			16'he6d6: y = 16'hfe01;
			16'he6d7: y = 16'hfe01;
			16'he6d8: y = 16'hfe01;
			16'he6d9: y = 16'hfe01;
			16'he6da: y = 16'hfe01;
			16'he6db: y = 16'hfe01;
			16'he6dc: y = 16'hfe01;
			16'he6dd: y = 16'hfe01;
			16'he6de: y = 16'hfe01;
			16'he6df: y = 16'hfe01;
			16'he6e0: y = 16'hfe01;
			16'he6e1: y = 16'hfe01;
			16'he6e2: y = 16'hfe01;
			16'he6e3: y = 16'hfe01;
			16'he6e4: y = 16'hfe01;
			16'he6e5: y = 16'hfe01;
			16'he6e6: y = 16'hfe01;
			16'he6e7: y = 16'hfe01;
			16'he6e8: y = 16'hfe01;
			16'he6e9: y = 16'hfe01;
			16'he6ea: y = 16'hfe01;
			16'he6eb: y = 16'hfe01;
			16'he6ec: y = 16'hfe01;
			16'he6ed: y = 16'hfe01;
			16'he6ee: y = 16'hfe01;
			16'he6ef: y = 16'hfe01;
			16'he6f0: y = 16'hfe01;
			16'he6f1: y = 16'hfe01;
			16'he6f2: y = 16'hfe01;
			16'he6f3: y = 16'hfe01;
			16'he6f4: y = 16'hfe01;
			16'he6f5: y = 16'hfe01;
			16'he6f6: y = 16'hfe01;
			16'he6f7: y = 16'hfe01;
			16'he6f8: y = 16'hfe01;
			16'he6f9: y = 16'hfe01;
			16'he6fa: y = 16'hfe01;
			16'he6fb: y = 16'hfe01;
			16'he6fc: y = 16'hfe01;
			16'he6fd: y = 16'hfe01;
			16'he6fe: y = 16'hfe01;
			16'he6ff: y = 16'hfe01;
			16'he700: y = 16'hfe01;
			16'he701: y = 16'hfe01;
			16'he702: y = 16'hfe01;
			16'he703: y = 16'hfe01;
			16'he704: y = 16'hfe01;
			16'he705: y = 16'hfe01;
			16'he706: y = 16'hfe01;
			16'he707: y = 16'hfe01;
			16'he708: y = 16'hfe01;
			16'he709: y = 16'hfe01;
			16'he70a: y = 16'hfe01;
			16'he70b: y = 16'hfe01;
			16'he70c: y = 16'hfe01;
			16'he70d: y = 16'hfe01;
			16'he70e: y = 16'hfe01;
			16'he70f: y = 16'hfe01;
			16'he710: y = 16'hfe01;
			16'he711: y = 16'hfe01;
			16'he712: y = 16'hfe01;
			16'he713: y = 16'hfe01;
			16'he714: y = 16'hfe01;
			16'he715: y = 16'hfe01;
			16'he716: y = 16'hfe01;
			16'he717: y = 16'hfe01;
			16'he718: y = 16'hfe01;
			16'he719: y = 16'hfe01;
			16'he71a: y = 16'hfe01;
			16'he71b: y = 16'hfe01;
			16'he71c: y = 16'hfe01;
			16'he71d: y = 16'hfe01;
			16'he71e: y = 16'hfe01;
			16'he71f: y = 16'hfe01;
			16'he720: y = 16'hfe01;
			16'he721: y = 16'hfe01;
			16'he722: y = 16'hfe01;
			16'he723: y = 16'hfe01;
			16'he724: y = 16'hfe01;
			16'he725: y = 16'hfe01;
			16'he726: y = 16'hfe01;
			16'he727: y = 16'hfe01;
			16'he728: y = 16'hfe01;
			16'he729: y = 16'hfe01;
			16'he72a: y = 16'hfe01;
			16'he72b: y = 16'hfe01;
			16'he72c: y = 16'hfe01;
			16'he72d: y = 16'hfe01;
			16'he72e: y = 16'hfe01;
			16'he72f: y = 16'hfe01;
			16'he730: y = 16'hfe01;
			16'he731: y = 16'hfe01;
			16'he732: y = 16'hfe01;
			16'he733: y = 16'hfe01;
			16'he734: y = 16'hfe01;
			16'he735: y = 16'hfe01;
			16'he736: y = 16'hfe01;
			16'he737: y = 16'hfe01;
			16'he738: y = 16'hfe01;
			16'he739: y = 16'hfe01;
			16'he73a: y = 16'hfe01;
			16'he73b: y = 16'hfe01;
			16'he73c: y = 16'hfe01;
			16'he73d: y = 16'hfe01;
			16'he73e: y = 16'hfe01;
			16'he73f: y = 16'hfe01;
			16'he740: y = 16'hfe01;
			16'he741: y = 16'hfe01;
			16'he742: y = 16'hfe01;
			16'he743: y = 16'hfe01;
			16'he744: y = 16'hfe01;
			16'he745: y = 16'hfe01;
			16'he746: y = 16'hfe01;
			16'he747: y = 16'hfe01;
			16'he748: y = 16'hfe01;
			16'he749: y = 16'hfe01;
			16'he74a: y = 16'hfe01;
			16'he74b: y = 16'hfe01;
			16'he74c: y = 16'hfe01;
			16'he74d: y = 16'hfe01;
			16'he74e: y = 16'hfe01;
			16'he74f: y = 16'hfe01;
			16'he750: y = 16'hfe01;
			16'he751: y = 16'hfe01;
			16'he752: y = 16'hfe01;
			16'he753: y = 16'hfe01;
			16'he754: y = 16'hfe01;
			16'he755: y = 16'hfe01;
			16'he756: y = 16'hfe01;
			16'he757: y = 16'hfe01;
			16'he758: y = 16'hfe01;
			16'he759: y = 16'hfe01;
			16'he75a: y = 16'hfe01;
			16'he75b: y = 16'hfe01;
			16'he75c: y = 16'hfe01;
			16'he75d: y = 16'hfe01;
			16'he75e: y = 16'hfe01;
			16'he75f: y = 16'hfe01;
			16'he760: y = 16'hfe01;
			16'he761: y = 16'hfe01;
			16'he762: y = 16'hfe01;
			16'he763: y = 16'hfe01;
			16'he764: y = 16'hfe01;
			16'he765: y = 16'hfe01;
			16'he766: y = 16'hfe01;
			16'he767: y = 16'hfe01;
			16'he768: y = 16'hfe01;
			16'he769: y = 16'hfe01;
			16'he76a: y = 16'hfe01;
			16'he76b: y = 16'hfe01;
			16'he76c: y = 16'hfe01;
			16'he76d: y = 16'hfe01;
			16'he76e: y = 16'hfe01;
			16'he76f: y = 16'hfe01;
			16'he770: y = 16'hfe01;
			16'he771: y = 16'hfe01;
			16'he772: y = 16'hfe01;
			16'he773: y = 16'hfe01;
			16'he774: y = 16'hfe01;
			16'he775: y = 16'hfe01;
			16'he776: y = 16'hfe01;
			16'he777: y = 16'hfe01;
			16'he778: y = 16'hfe01;
			16'he779: y = 16'hfe01;
			16'he77a: y = 16'hfe01;
			16'he77b: y = 16'hfe01;
			16'he77c: y = 16'hfe01;
			16'he77d: y = 16'hfe01;
			16'he77e: y = 16'hfe01;
			16'he77f: y = 16'hfe01;
			16'he780: y = 16'hfe01;
			16'he781: y = 16'hfe01;
			16'he782: y = 16'hfe01;
			16'he783: y = 16'hfe01;
			16'he784: y = 16'hfe01;
			16'he785: y = 16'hfe01;
			16'he786: y = 16'hfe01;
			16'he787: y = 16'hfe01;
			16'he788: y = 16'hfe01;
			16'he789: y = 16'hfe01;
			16'he78a: y = 16'hfe01;
			16'he78b: y = 16'hfe01;
			16'he78c: y = 16'hfe01;
			16'he78d: y = 16'hfe01;
			16'he78e: y = 16'hfe01;
			16'he78f: y = 16'hfe01;
			16'he790: y = 16'hfe01;
			16'he791: y = 16'hfe01;
			16'he792: y = 16'hfe01;
			16'he793: y = 16'hfe01;
			16'he794: y = 16'hfe01;
			16'he795: y = 16'hfe01;
			16'he796: y = 16'hfe01;
			16'he797: y = 16'hfe01;
			16'he798: y = 16'hfe01;
			16'he799: y = 16'hfe01;
			16'he79a: y = 16'hfe01;
			16'he79b: y = 16'hfe01;
			16'he79c: y = 16'hfe01;
			16'he79d: y = 16'hfe01;
			16'he79e: y = 16'hfe01;
			16'he79f: y = 16'hfe01;
			16'he7a0: y = 16'hfe01;
			16'he7a1: y = 16'hfe01;
			16'he7a2: y = 16'hfe01;
			16'he7a3: y = 16'hfe01;
			16'he7a4: y = 16'hfe01;
			16'he7a5: y = 16'hfe01;
			16'he7a6: y = 16'hfe01;
			16'he7a7: y = 16'hfe01;
			16'he7a8: y = 16'hfe01;
			16'he7a9: y = 16'hfe01;
			16'he7aa: y = 16'hfe01;
			16'he7ab: y = 16'hfe01;
			16'he7ac: y = 16'hfe01;
			16'he7ad: y = 16'hfe01;
			16'he7ae: y = 16'hfe01;
			16'he7af: y = 16'hfe01;
			16'he7b0: y = 16'hfe01;
			16'he7b1: y = 16'hfe01;
			16'he7b2: y = 16'hfe01;
			16'he7b3: y = 16'hfe01;
			16'he7b4: y = 16'hfe01;
			16'he7b5: y = 16'hfe01;
			16'he7b6: y = 16'hfe01;
			16'he7b7: y = 16'hfe01;
			16'he7b8: y = 16'hfe01;
			16'he7b9: y = 16'hfe01;
			16'he7ba: y = 16'hfe01;
			16'he7bb: y = 16'hfe01;
			16'he7bc: y = 16'hfe01;
			16'he7bd: y = 16'hfe01;
			16'he7be: y = 16'hfe01;
			16'he7bf: y = 16'hfe01;
			16'he7c0: y = 16'hfe01;
			16'he7c1: y = 16'hfe01;
			16'he7c2: y = 16'hfe01;
			16'he7c3: y = 16'hfe01;
			16'he7c4: y = 16'hfe01;
			16'he7c5: y = 16'hfe01;
			16'he7c6: y = 16'hfe01;
			16'he7c7: y = 16'hfe01;
			16'he7c8: y = 16'hfe01;
			16'he7c9: y = 16'hfe01;
			16'he7ca: y = 16'hfe01;
			16'he7cb: y = 16'hfe01;
			16'he7cc: y = 16'hfe01;
			16'he7cd: y = 16'hfe01;
			16'he7ce: y = 16'hfe01;
			16'he7cf: y = 16'hfe01;
			16'he7d0: y = 16'hfe01;
			16'he7d1: y = 16'hfe01;
			16'he7d2: y = 16'hfe01;
			16'he7d3: y = 16'hfe01;
			16'he7d4: y = 16'hfe01;
			16'he7d5: y = 16'hfe01;
			16'he7d6: y = 16'hfe01;
			16'he7d7: y = 16'hfe01;
			16'he7d8: y = 16'hfe01;
			16'he7d9: y = 16'hfe01;
			16'he7da: y = 16'hfe01;
			16'he7db: y = 16'hfe01;
			16'he7dc: y = 16'hfe01;
			16'he7dd: y = 16'hfe01;
			16'he7de: y = 16'hfe01;
			16'he7df: y = 16'hfe01;
			16'he7e0: y = 16'hfe01;
			16'he7e1: y = 16'hfe01;
			16'he7e2: y = 16'hfe01;
			16'he7e3: y = 16'hfe01;
			16'he7e4: y = 16'hfe01;
			16'he7e5: y = 16'hfe01;
			16'he7e6: y = 16'hfe01;
			16'he7e7: y = 16'hfe01;
			16'he7e8: y = 16'hfe01;
			16'he7e9: y = 16'hfe01;
			16'he7ea: y = 16'hfe01;
			16'he7eb: y = 16'hfe01;
			16'he7ec: y = 16'hfe01;
			16'he7ed: y = 16'hfe01;
			16'he7ee: y = 16'hfe01;
			16'he7ef: y = 16'hfe01;
			16'he7f0: y = 16'hfe01;
			16'he7f1: y = 16'hfe01;
			16'he7f2: y = 16'hfe01;
			16'he7f3: y = 16'hfe01;
			16'he7f4: y = 16'hfe01;
			16'he7f5: y = 16'hfe01;
			16'he7f6: y = 16'hfe01;
			16'he7f7: y = 16'hfe01;
			16'he7f8: y = 16'hfe01;
			16'he7f9: y = 16'hfe01;
			16'he7fa: y = 16'hfe01;
			16'he7fb: y = 16'hfe01;
			16'he7fc: y = 16'hfe01;
			16'he7fd: y = 16'hfe01;
			16'he7fe: y = 16'hfe01;
			16'he7ff: y = 16'hfe01;
			16'he800: y = 16'hfe01;
			16'he801: y = 16'hfe01;
			16'he802: y = 16'hfe01;
			16'he803: y = 16'hfe01;
			16'he804: y = 16'hfe01;
			16'he805: y = 16'hfe01;
			16'he806: y = 16'hfe01;
			16'he807: y = 16'hfe01;
			16'he808: y = 16'hfe01;
			16'he809: y = 16'hfe01;
			16'he80a: y = 16'hfe01;
			16'he80b: y = 16'hfe01;
			16'he80c: y = 16'hfe01;
			16'he80d: y = 16'hfe01;
			16'he80e: y = 16'hfe01;
			16'he80f: y = 16'hfe01;
			16'he810: y = 16'hfe01;
			16'he811: y = 16'hfe01;
			16'he812: y = 16'hfe01;
			16'he813: y = 16'hfe01;
			16'he814: y = 16'hfe01;
			16'he815: y = 16'hfe01;
			16'he816: y = 16'hfe01;
			16'he817: y = 16'hfe01;
			16'he818: y = 16'hfe01;
			16'he819: y = 16'hfe01;
			16'he81a: y = 16'hfe01;
			16'he81b: y = 16'hfe01;
			16'he81c: y = 16'hfe01;
			16'he81d: y = 16'hfe01;
			16'he81e: y = 16'hfe01;
			16'he81f: y = 16'hfe01;
			16'he820: y = 16'hfe01;
			16'he821: y = 16'hfe01;
			16'he822: y = 16'hfe01;
			16'he823: y = 16'hfe01;
			16'he824: y = 16'hfe01;
			16'he825: y = 16'hfe01;
			16'he826: y = 16'hfe01;
			16'he827: y = 16'hfe01;
			16'he828: y = 16'hfe01;
			16'he829: y = 16'hfe01;
			16'he82a: y = 16'hfe01;
			16'he82b: y = 16'hfe01;
			16'he82c: y = 16'hfe01;
			16'he82d: y = 16'hfe01;
			16'he82e: y = 16'hfe01;
			16'he82f: y = 16'hfe01;
			16'he830: y = 16'hfe01;
			16'he831: y = 16'hfe01;
			16'he832: y = 16'hfe01;
			16'he833: y = 16'hfe01;
			16'he834: y = 16'hfe01;
			16'he835: y = 16'hfe01;
			16'he836: y = 16'hfe01;
			16'he837: y = 16'hfe01;
			16'he838: y = 16'hfe01;
			16'he839: y = 16'hfe01;
			16'he83a: y = 16'hfe01;
			16'he83b: y = 16'hfe01;
			16'he83c: y = 16'hfe01;
			16'he83d: y = 16'hfe01;
			16'he83e: y = 16'hfe01;
			16'he83f: y = 16'hfe01;
			16'he840: y = 16'hfe01;
			16'he841: y = 16'hfe01;
			16'he842: y = 16'hfe01;
			16'he843: y = 16'hfe01;
			16'he844: y = 16'hfe01;
			16'he845: y = 16'hfe01;
			16'he846: y = 16'hfe01;
			16'he847: y = 16'hfe01;
			16'he848: y = 16'hfe01;
			16'he849: y = 16'hfe01;
			16'he84a: y = 16'hfe01;
			16'he84b: y = 16'hfe01;
			16'he84c: y = 16'hfe01;
			16'he84d: y = 16'hfe01;
			16'he84e: y = 16'hfe01;
			16'he84f: y = 16'hfe01;
			16'he850: y = 16'hfe01;
			16'he851: y = 16'hfe01;
			16'he852: y = 16'hfe01;
			16'he853: y = 16'hfe01;
			16'he854: y = 16'hfe01;
			16'he855: y = 16'hfe01;
			16'he856: y = 16'hfe01;
			16'he857: y = 16'hfe01;
			16'he858: y = 16'hfe01;
			16'he859: y = 16'hfe01;
			16'he85a: y = 16'hfe01;
			16'he85b: y = 16'hfe01;
			16'he85c: y = 16'hfe01;
			16'he85d: y = 16'hfe01;
			16'he85e: y = 16'hfe01;
			16'he85f: y = 16'hfe01;
			16'he860: y = 16'hfe01;
			16'he861: y = 16'hfe01;
			16'he862: y = 16'hfe01;
			16'he863: y = 16'hfe01;
			16'he864: y = 16'hfe01;
			16'he865: y = 16'hfe01;
			16'he866: y = 16'hfe01;
			16'he867: y = 16'hfe01;
			16'he868: y = 16'hfe01;
			16'he869: y = 16'hfe01;
			16'he86a: y = 16'hfe01;
			16'he86b: y = 16'hfe01;
			16'he86c: y = 16'hfe01;
			16'he86d: y = 16'hfe01;
			16'he86e: y = 16'hfe01;
			16'he86f: y = 16'hfe01;
			16'he870: y = 16'hfe01;
			16'he871: y = 16'hfe01;
			16'he872: y = 16'hfe01;
			16'he873: y = 16'hfe01;
			16'he874: y = 16'hfe01;
			16'he875: y = 16'hfe01;
			16'he876: y = 16'hfe01;
			16'he877: y = 16'hfe01;
			16'he878: y = 16'hfe01;
			16'he879: y = 16'hfe01;
			16'he87a: y = 16'hfe01;
			16'he87b: y = 16'hfe01;
			16'he87c: y = 16'hfe01;
			16'he87d: y = 16'hfe01;
			16'he87e: y = 16'hfe01;
			16'he87f: y = 16'hfe01;
			16'he880: y = 16'hfe01;
			16'he881: y = 16'hfe01;
			16'he882: y = 16'hfe01;
			16'he883: y = 16'hfe01;
			16'he884: y = 16'hfe01;
			16'he885: y = 16'hfe01;
			16'he886: y = 16'hfe01;
			16'he887: y = 16'hfe01;
			16'he888: y = 16'hfe01;
			16'he889: y = 16'hfe01;
			16'he88a: y = 16'hfe01;
			16'he88b: y = 16'hfe01;
			16'he88c: y = 16'hfe01;
			16'he88d: y = 16'hfe01;
			16'he88e: y = 16'hfe01;
			16'he88f: y = 16'hfe01;
			16'he890: y = 16'hfe01;
			16'he891: y = 16'hfe01;
			16'he892: y = 16'hfe01;
			16'he893: y = 16'hfe01;
			16'he894: y = 16'hfe01;
			16'he895: y = 16'hfe01;
			16'he896: y = 16'hfe01;
			16'he897: y = 16'hfe01;
			16'he898: y = 16'hfe01;
			16'he899: y = 16'hfe01;
			16'he89a: y = 16'hfe01;
			16'he89b: y = 16'hfe01;
			16'he89c: y = 16'hfe01;
			16'he89d: y = 16'hfe01;
			16'he89e: y = 16'hfe01;
			16'he89f: y = 16'hfe01;
			16'he8a0: y = 16'hfe01;
			16'he8a1: y = 16'hfe01;
			16'he8a2: y = 16'hfe01;
			16'he8a3: y = 16'hfe01;
			16'he8a4: y = 16'hfe01;
			16'he8a5: y = 16'hfe01;
			16'he8a6: y = 16'hfe01;
			16'he8a7: y = 16'hfe01;
			16'he8a8: y = 16'hfe01;
			16'he8a9: y = 16'hfe01;
			16'he8aa: y = 16'hfe01;
			16'he8ab: y = 16'hfe01;
			16'he8ac: y = 16'hfe01;
			16'he8ad: y = 16'hfe01;
			16'he8ae: y = 16'hfe01;
			16'he8af: y = 16'hfe01;
			16'he8b0: y = 16'hfe01;
			16'he8b1: y = 16'hfe01;
			16'he8b2: y = 16'hfe01;
			16'he8b3: y = 16'hfe01;
			16'he8b4: y = 16'hfe01;
			16'he8b5: y = 16'hfe01;
			16'he8b6: y = 16'hfe01;
			16'he8b7: y = 16'hfe01;
			16'he8b8: y = 16'hfe01;
			16'he8b9: y = 16'hfe01;
			16'he8ba: y = 16'hfe01;
			16'he8bb: y = 16'hfe01;
			16'he8bc: y = 16'hfe01;
			16'he8bd: y = 16'hfe01;
			16'he8be: y = 16'hfe01;
			16'he8bf: y = 16'hfe01;
			16'he8c0: y = 16'hfe01;
			16'he8c1: y = 16'hfe01;
			16'he8c2: y = 16'hfe01;
			16'he8c3: y = 16'hfe01;
			16'he8c4: y = 16'hfe01;
			16'he8c5: y = 16'hfe01;
			16'he8c6: y = 16'hfe01;
			16'he8c7: y = 16'hfe01;
			16'he8c8: y = 16'hfe01;
			16'he8c9: y = 16'hfe01;
			16'he8ca: y = 16'hfe01;
			16'he8cb: y = 16'hfe01;
			16'he8cc: y = 16'hfe01;
			16'he8cd: y = 16'hfe01;
			16'he8ce: y = 16'hfe01;
			16'he8cf: y = 16'hfe01;
			16'he8d0: y = 16'hfe01;
			16'he8d1: y = 16'hfe01;
			16'he8d2: y = 16'hfe01;
			16'he8d3: y = 16'hfe01;
			16'he8d4: y = 16'hfe01;
			16'he8d5: y = 16'hfe01;
			16'he8d6: y = 16'hfe01;
			16'he8d7: y = 16'hfe01;
			16'he8d8: y = 16'hfe01;
			16'he8d9: y = 16'hfe01;
			16'he8da: y = 16'hfe01;
			16'he8db: y = 16'hfe01;
			16'he8dc: y = 16'hfe01;
			16'he8dd: y = 16'hfe01;
			16'he8de: y = 16'hfe01;
			16'he8df: y = 16'hfe01;
			16'he8e0: y = 16'hfe01;
			16'he8e1: y = 16'hfe01;
			16'he8e2: y = 16'hfe01;
			16'he8e3: y = 16'hfe01;
			16'he8e4: y = 16'hfe01;
			16'he8e5: y = 16'hfe01;
			16'he8e6: y = 16'hfe01;
			16'he8e7: y = 16'hfe01;
			16'he8e8: y = 16'hfe01;
			16'he8e9: y = 16'hfe01;
			16'he8ea: y = 16'hfe01;
			16'he8eb: y = 16'hfe01;
			16'he8ec: y = 16'hfe01;
			16'he8ed: y = 16'hfe01;
			16'he8ee: y = 16'hfe01;
			16'he8ef: y = 16'hfe01;
			16'he8f0: y = 16'hfe01;
			16'he8f1: y = 16'hfe01;
			16'he8f2: y = 16'hfe01;
			16'he8f3: y = 16'hfe01;
			16'he8f4: y = 16'hfe01;
			16'he8f5: y = 16'hfe01;
			16'he8f6: y = 16'hfe01;
			16'he8f7: y = 16'hfe01;
			16'he8f8: y = 16'hfe01;
			16'he8f9: y = 16'hfe01;
			16'he8fa: y = 16'hfe01;
			16'he8fb: y = 16'hfe01;
			16'he8fc: y = 16'hfe01;
			16'he8fd: y = 16'hfe01;
			16'he8fe: y = 16'hfe01;
			16'he8ff: y = 16'hfe01;
			16'he900: y = 16'hfe01;
			16'he901: y = 16'hfe01;
			16'he902: y = 16'hfe01;
			16'he903: y = 16'hfe01;
			16'he904: y = 16'hfe01;
			16'he905: y = 16'hfe01;
			16'he906: y = 16'hfe01;
			16'he907: y = 16'hfe01;
			16'he908: y = 16'hfe01;
			16'he909: y = 16'hfe01;
			16'he90a: y = 16'hfe01;
			16'he90b: y = 16'hfe01;
			16'he90c: y = 16'hfe01;
			16'he90d: y = 16'hfe01;
			16'he90e: y = 16'hfe01;
			16'he90f: y = 16'hfe01;
			16'he910: y = 16'hfe01;
			16'he911: y = 16'hfe01;
			16'he912: y = 16'hfe01;
			16'he913: y = 16'hfe01;
			16'he914: y = 16'hfe01;
			16'he915: y = 16'hfe01;
			16'he916: y = 16'hfe01;
			16'he917: y = 16'hfe01;
			16'he918: y = 16'hfe01;
			16'he919: y = 16'hfe01;
			16'he91a: y = 16'hfe01;
			16'he91b: y = 16'hfe01;
			16'he91c: y = 16'hfe01;
			16'he91d: y = 16'hfe01;
			16'he91e: y = 16'hfe01;
			16'he91f: y = 16'hfe01;
			16'he920: y = 16'hfe01;
			16'he921: y = 16'hfe01;
			16'he922: y = 16'hfe01;
			16'he923: y = 16'hfe01;
			16'he924: y = 16'hfe01;
			16'he925: y = 16'hfe01;
			16'he926: y = 16'hfe01;
			16'he927: y = 16'hfe01;
			16'he928: y = 16'hfe01;
			16'he929: y = 16'hfe01;
			16'he92a: y = 16'hfe01;
			16'he92b: y = 16'hfe01;
			16'he92c: y = 16'hfe01;
			16'he92d: y = 16'hfe01;
			16'he92e: y = 16'hfe01;
			16'he92f: y = 16'hfe01;
			16'he930: y = 16'hfe01;
			16'he931: y = 16'hfe01;
			16'he932: y = 16'hfe01;
			16'he933: y = 16'hfe01;
			16'he934: y = 16'hfe01;
			16'he935: y = 16'hfe01;
			16'he936: y = 16'hfe01;
			16'he937: y = 16'hfe01;
			16'he938: y = 16'hfe01;
			16'he939: y = 16'hfe01;
			16'he93a: y = 16'hfe01;
			16'he93b: y = 16'hfe01;
			16'he93c: y = 16'hfe01;
			16'he93d: y = 16'hfe01;
			16'he93e: y = 16'hfe01;
			16'he93f: y = 16'hfe01;
			16'he940: y = 16'hfe01;
			16'he941: y = 16'hfe01;
			16'he942: y = 16'hfe01;
			16'he943: y = 16'hfe01;
			16'he944: y = 16'hfe01;
			16'he945: y = 16'hfe01;
			16'he946: y = 16'hfe01;
			16'he947: y = 16'hfe01;
			16'he948: y = 16'hfe01;
			16'he949: y = 16'hfe01;
			16'he94a: y = 16'hfe01;
			16'he94b: y = 16'hfe01;
			16'he94c: y = 16'hfe01;
			16'he94d: y = 16'hfe01;
			16'he94e: y = 16'hfe01;
			16'he94f: y = 16'hfe01;
			16'he950: y = 16'hfe01;
			16'he951: y = 16'hfe01;
			16'he952: y = 16'hfe01;
			16'he953: y = 16'hfe01;
			16'he954: y = 16'hfe01;
			16'he955: y = 16'hfe01;
			16'he956: y = 16'hfe01;
			16'he957: y = 16'hfe01;
			16'he958: y = 16'hfe01;
			16'he959: y = 16'hfe01;
			16'he95a: y = 16'hfe01;
			16'he95b: y = 16'hfe01;
			16'he95c: y = 16'hfe01;
			16'he95d: y = 16'hfe01;
			16'he95e: y = 16'hfe01;
			16'he95f: y = 16'hfe01;
			16'he960: y = 16'hfe01;
			16'he961: y = 16'hfe01;
			16'he962: y = 16'hfe01;
			16'he963: y = 16'hfe01;
			16'he964: y = 16'hfe01;
			16'he965: y = 16'hfe01;
			16'he966: y = 16'hfe01;
			16'he967: y = 16'hfe01;
			16'he968: y = 16'hfe01;
			16'he969: y = 16'hfe01;
			16'he96a: y = 16'hfe01;
			16'he96b: y = 16'hfe01;
			16'he96c: y = 16'hfe01;
			16'he96d: y = 16'hfe01;
			16'he96e: y = 16'hfe01;
			16'he96f: y = 16'hfe01;
			16'he970: y = 16'hfe01;
			16'he971: y = 16'hfe01;
			16'he972: y = 16'hfe01;
			16'he973: y = 16'hfe01;
			16'he974: y = 16'hfe01;
			16'he975: y = 16'hfe01;
			16'he976: y = 16'hfe01;
			16'he977: y = 16'hfe01;
			16'he978: y = 16'hfe01;
			16'he979: y = 16'hfe01;
			16'he97a: y = 16'hfe01;
			16'he97b: y = 16'hfe01;
			16'he97c: y = 16'hfe01;
			16'he97d: y = 16'hfe01;
			16'he97e: y = 16'hfe01;
			16'he97f: y = 16'hfe01;
			16'he980: y = 16'hfe01;
			16'he981: y = 16'hfe01;
			16'he982: y = 16'hfe01;
			16'he983: y = 16'hfe01;
			16'he984: y = 16'hfe01;
			16'he985: y = 16'hfe01;
			16'he986: y = 16'hfe01;
			16'he987: y = 16'hfe01;
			16'he988: y = 16'hfe01;
			16'he989: y = 16'hfe01;
			16'he98a: y = 16'hfe01;
			16'he98b: y = 16'hfe01;
			16'he98c: y = 16'hfe01;
			16'he98d: y = 16'hfe01;
			16'he98e: y = 16'hfe01;
			16'he98f: y = 16'hfe01;
			16'he990: y = 16'hfe01;
			16'he991: y = 16'hfe01;
			16'he992: y = 16'hfe01;
			16'he993: y = 16'hfe01;
			16'he994: y = 16'hfe01;
			16'he995: y = 16'hfe01;
			16'he996: y = 16'hfe01;
			16'he997: y = 16'hfe01;
			16'he998: y = 16'hfe01;
			16'he999: y = 16'hfe01;
			16'he99a: y = 16'hfe01;
			16'he99b: y = 16'hfe01;
			16'he99c: y = 16'hfe01;
			16'he99d: y = 16'hfe01;
			16'he99e: y = 16'hfe01;
			16'he99f: y = 16'hfe01;
			16'he9a0: y = 16'hfe01;
			16'he9a1: y = 16'hfe01;
			16'he9a2: y = 16'hfe01;
			16'he9a3: y = 16'hfe01;
			16'he9a4: y = 16'hfe01;
			16'he9a5: y = 16'hfe01;
			16'he9a6: y = 16'hfe01;
			16'he9a7: y = 16'hfe01;
			16'he9a8: y = 16'hfe01;
			16'he9a9: y = 16'hfe01;
			16'he9aa: y = 16'hfe01;
			16'he9ab: y = 16'hfe01;
			16'he9ac: y = 16'hfe01;
			16'he9ad: y = 16'hfe01;
			16'he9ae: y = 16'hfe01;
			16'he9af: y = 16'hfe01;
			16'he9b0: y = 16'hfe01;
			16'he9b1: y = 16'hfe01;
			16'he9b2: y = 16'hfe01;
			16'he9b3: y = 16'hfe01;
			16'he9b4: y = 16'hfe01;
			16'he9b5: y = 16'hfe01;
			16'he9b6: y = 16'hfe01;
			16'he9b7: y = 16'hfe01;
			16'he9b8: y = 16'hfe01;
			16'he9b9: y = 16'hfe01;
			16'he9ba: y = 16'hfe01;
			16'he9bb: y = 16'hfe01;
			16'he9bc: y = 16'hfe01;
			16'he9bd: y = 16'hfe01;
			16'he9be: y = 16'hfe01;
			16'he9bf: y = 16'hfe01;
			16'he9c0: y = 16'hfe01;
			16'he9c1: y = 16'hfe01;
			16'he9c2: y = 16'hfe01;
			16'he9c3: y = 16'hfe01;
			16'he9c4: y = 16'hfe01;
			16'he9c5: y = 16'hfe01;
			16'he9c6: y = 16'hfe01;
			16'he9c7: y = 16'hfe01;
			16'he9c8: y = 16'hfe01;
			16'he9c9: y = 16'hfe01;
			16'he9ca: y = 16'hfe01;
			16'he9cb: y = 16'hfe01;
			16'he9cc: y = 16'hfe01;
			16'he9cd: y = 16'hfe01;
			16'he9ce: y = 16'hfe01;
			16'he9cf: y = 16'hfe01;
			16'he9d0: y = 16'hfe01;
			16'he9d1: y = 16'hfe01;
			16'he9d2: y = 16'hfe01;
			16'he9d3: y = 16'hfe01;
			16'he9d4: y = 16'hfe01;
			16'he9d5: y = 16'hfe01;
			16'he9d6: y = 16'hfe01;
			16'he9d7: y = 16'hfe01;
			16'he9d8: y = 16'hfe01;
			16'he9d9: y = 16'hfe01;
			16'he9da: y = 16'hfe01;
			16'he9db: y = 16'hfe01;
			16'he9dc: y = 16'hfe01;
			16'he9dd: y = 16'hfe01;
			16'he9de: y = 16'hfe01;
			16'he9df: y = 16'hfe01;
			16'he9e0: y = 16'hfe01;
			16'he9e1: y = 16'hfe01;
			16'he9e2: y = 16'hfe01;
			16'he9e3: y = 16'hfe01;
			16'he9e4: y = 16'hfe01;
			16'he9e5: y = 16'hfe01;
			16'he9e6: y = 16'hfe01;
			16'he9e7: y = 16'hfe01;
			16'he9e8: y = 16'hfe01;
			16'he9e9: y = 16'hfe01;
			16'he9ea: y = 16'hfe01;
			16'he9eb: y = 16'hfe01;
			16'he9ec: y = 16'hfe01;
			16'he9ed: y = 16'hfe01;
			16'he9ee: y = 16'hfe01;
			16'he9ef: y = 16'hfe01;
			16'he9f0: y = 16'hfe01;
			16'he9f1: y = 16'hfe01;
			16'he9f2: y = 16'hfe01;
			16'he9f3: y = 16'hfe01;
			16'he9f4: y = 16'hfe01;
			16'he9f5: y = 16'hfe01;
			16'he9f6: y = 16'hfe01;
			16'he9f7: y = 16'hfe01;
			16'he9f8: y = 16'hfe01;
			16'he9f9: y = 16'hfe01;
			16'he9fa: y = 16'hfe01;
			16'he9fb: y = 16'hfe01;
			16'he9fc: y = 16'hfe01;
			16'he9fd: y = 16'hfe01;
			16'he9fe: y = 16'hfe01;
			16'he9ff: y = 16'hfe01;
			16'hea00: y = 16'hfe01;
			16'hea01: y = 16'hfe01;
			16'hea02: y = 16'hfe01;
			16'hea03: y = 16'hfe01;
			16'hea04: y = 16'hfe01;
			16'hea05: y = 16'hfe01;
			16'hea06: y = 16'hfe01;
			16'hea07: y = 16'hfe01;
			16'hea08: y = 16'hfe01;
			16'hea09: y = 16'hfe01;
			16'hea0a: y = 16'hfe01;
			16'hea0b: y = 16'hfe01;
			16'hea0c: y = 16'hfe01;
			16'hea0d: y = 16'hfe01;
			16'hea0e: y = 16'hfe01;
			16'hea0f: y = 16'hfe01;
			16'hea10: y = 16'hfe01;
			16'hea11: y = 16'hfe01;
			16'hea12: y = 16'hfe01;
			16'hea13: y = 16'hfe01;
			16'hea14: y = 16'hfe01;
			16'hea15: y = 16'hfe01;
			16'hea16: y = 16'hfe01;
			16'hea17: y = 16'hfe01;
			16'hea18: y = 16'hfe01;
			16'hea19: y = 16'hfe01;
			16'hea1a: y = 16'hfe01;
			16'hea1b: y = 16'hfe01;
			16'hea1c: y = 16'hfe01;
			16'hea1d: y = 16'hfe01;
			16'hea1e: y = 16'hfe01;
			16'hea1f: y = 16'hfe01;
			16'hea20: y = 16'hfe01;
			16'hea21: y = 16'hfe01;
			16'hea22: y = 16'hfe01;
			16'hea23: y = 16'hfe01;
			16'hea24: y = 16'hfe01;
			16'hea25: y = 16'hfe01;
			16'hea26: y = 16'hfe01;
			16'hea27: y = 16'hfe01;
			16'hea28: y = 16'hfe01;
			16'hea29: y = 16'hfe01;
			16'hea2a: y = 16'hfe01;
			16'hea2b: y = 16'hfe01;
			16'hea2c: y = 16'hfe01;
			16'hea2d: y = 16'hfe01;
			16'hea2e: y = 16'hfe01;
			16'hea2f: y = 16'hfe01;
			16'hea30: y = 16'hfe01;
			16'hea31: y = 16'hfe01;
			16'hea32: y = 16'hfe01;
			16'hea33: y = 16'hfe01;
			16'hea34: y = 16'hfe01;
			16'hea35: y = 16'hfe01;
			16'hea36: y = 16'hfe01;
			16'hea37: y = 16'hfe01;
			16'hea38: y = 16'hfe01;
			16'hea39: y = 16'hfe01;
			16'hea3a: y = 16'hfe01;
			16'hea3b: y = 16'hfe01;
			16'hea3c: y = 16'hfe01;
			16'hea3d: y = 16'hfe01;
			16'hea3e: y = 16'hfe01;
			16'hea3f: y = 16'hfe01;
			16'hea40: y = 16'hfe01;
			16'hea41: y = 16'hfe01;
			16'hea42: y = 16'hfe01;
			16'hea43: y = 16'hfe01;
			16'hea44: y = 16'hfe01;
			16'hea45: y = 16'hfe01;
			16'hea46: y = 16'hfe01;
			16'hea47: y = 16'hfe01;
			16'hea48: y = 16'hfe01;
			16'hea49: y = 16'hfe01;
			16'hea4a: y = 16'hfe01;
			16'hea4b: y = 16'hfe01;
			16'hea4c: y = 16'hfe01;
			16'hea4d: y = 16'hfe01;
			16'hea4e: y = 16'hfe01;
			16'hea4f: y = 16'hfe01;
			16'hea50: y = 16'hfe01;
			16'hea51: y = 16'hfe01;
			16'hea52: y = 16'hfe01;
			16'hea53: y = 16'hfe01;
			16'hea54: y = 16'hfe01;
			16'hea55: y = 16'hfe01;
			16'hea56: y = 16'hfe01;
			16'hea57: y = 16'hfe01;
			16'hea58: y = 16'hfe01;
			16'hea59: y = 16'hfe01;
			16'hea5a: y = 16'hfe01;
			16'hea5b: y = 16'hfe01;
			16'hea5c: y = 16'hfe01;
			16'hea5d: y = 16'hfe01;
			16'hea5e: y = 16'hfe01;
			16'hea5f: y = 16'hfe01;
			16'hea60: y = 16'hfe01;
			16'hea61: y = 16'hfe01;
			16'hea62: y = 16'hfe01;
			16'hea63: y = 16'hfe01;
			16'hea64: y = 16'hfe01;
			16'hea65: y = 16'hfe01;
			16'hea66: y = 16'hfe01;
			16'hea67: y = 16'hfe01;
			16'hea68: y = 16'hfe01;
			16'hea69: y = 16'hfe01;
			16'hea6a: y = 16'hfe01;
			16'hea6b: y = 16'hfe01;
			16'hea6c: y = 16'hfe01;
			16'hea6d: y = 16'hfe01;
			16'hea6e: y = 16'hfe01;
			16'hea6f: y = 16'hfe01;
			16'hea70: y = 16'hfe01;
			16'hea71: y = 16'hfe01;
			16'hea72: y = 16'hfe01;
			16'hea73: y = 16'hfe01;
			16'hea74: y = 16'hfe01;
			16'hea75: y = 16'hfe01;
			16'hea76: y = 16'hfe01;
			16'hea77: y = 16'hfe01;
			16'hea78: y = 16'hfe01;
			16'hea79: y = 16'hfe01;
			16'hea7a: y = 16'hfe01;
			16'hea7b: y = 16'hfe01;
			16'hea7c: y = 16'hfe01;
			16'hea7d: y = 16'hfe01;
			16'hea7e: y = 16'hfe01;
			16'hea7f: y = 16'hfe01;
			16'hea80: y = 16'hfe01;
			16'hea81: y = 16'hfe01;
			16'hea82: y = 16'hfe01;
			16'hea83: y = 16'hfe01;
			16'hea84: y = 16'hfe01;
			16'hea85: y = 16'hfe01;
			16'hea86: y = 16'hfe01;
			16'hea87: y = 16'hfe01;
			16'hea88: y = 16'hfe01;
			16'hea89: y = 16'hfe01;
			16'hea8a: y = 16'hfe01;
			16'hea8b: y = 16'hfe01;
			16'hea8c: y = 16'hfe01;
			16'hea8d: y = 16'hfe01;
			16'hea8e: y = 16'hfe01;
			16'hea8f: y = 16'hfe01;
			16'hea90: y = 16'hfe01;
			16'hea91: y = 16'hfe01;
			16'hea92: y = 16'hfe01;
			16'hea93: y = 16'hfe01;
			16'hea94: y = 16'hfe01;
			16'hea95: y = 16'hfe01;
			16'hea96: y = 16'hfe01;
			16'hea97: y = 16'hfe01;
			16'hea98: y = 16'hfe01;
			16'hea99: y = 16'hfe01;
			16'hea9a: y = 16'hfe01;
			16'hea9b: y = 16'hfe01;
			16'hea9c: y = 16'hfe01;
			16'hea9d: y = 16'hfe01;
			16'hea9e: y = 16'hfe01;
			16'hea9f: y = 16'hfe01;
			16'heaa0: y = 16'hfe01;
			16'heaa1: y = 16'hfe01;
			16'heaa2: y = 16'hfe01;
			16'heaa3: y = 16'hfe01;
			16'heaa4: y = 16'hfe01;
			16'heaa5: y = 16'hfe01;
			16'heaa6: y = 16'hfe01;
			16'heaa7: y = 16'hfe01;
			16'heaa8: y = 16'hfe01;
			16'heaa9: y = 16'hfe01;
			16'heaaa: y = 16'hfe01;
			16'heaab: y = 16'hfe01;
			16'heaac: y = 16'hfe01;
			16'heaad: y = 16'hfe01;
			16'heaae: y = 16'hfe01;
			16'heaaf: y = 16'hfe01;
			16'heab0: y = 16'hfe01;
			16'heab1: y = 16'hfe01;
			16'heab2: y = 16'hfe01;
			16'heab3: y = 16'hfe01;
			16'heab4: y = 16'hfe01;
			16'heab5: y = 16'hfe01;
			16'heab6: y = 16'hfe01;
			16'heab7: y = 16'hfe01;
			16'heab8: y = 16'hfe01;
			16'heab9: y = 16'hfe01;
			16'heaba: y = 16'hfe01;
			16'heabb: y = 16'hfe01;
			16'heabc: y = 16'hfe01;
			16'heabd: y = 16'hfe01;
			16'heabe: y = 16'hfe01;
			16'heabf: y = 16'hfe01;
			16'heac0: y = 16'hfe01;
			16'heac1: y = 16'hfe01;
			16'heac2: y = 16'hfe01;
			16'heac3: y = 16'hfe01;
			16'heac4: y = 16'hfe01;
			16'heac5: y = 16'hfe01;
			16'heac6: y = 16'hfe01;
			16'heac7: y = 16'hfe01;
			16'heac8: y = 16'hfe01;
			16'heac9: y = 16'hfe01;
			16'heaca: y = 16'hfe01;
			16'heacb: y = 16'hfe01;
			16'heacc: y = 16'hfe01;
			16'heacd: y = 16'hfe01;
			16'heace: y = 16'hfe01;
			16'heacf: y = 16'hfe01;
			16'head0: y = 16'hfe01;
			16'head1: y = 16'hfe01;
			16'head2: y = 16'hfe01;
			16'head3: y = 16'hfe01;
			16'head4: y = 16'hfe01;
			16'head5: y = 16'hfe01;
			16'head6: y = 16'hfe01;
			16'head7: y = 16'hfe01;
			16'head8: y = 16'hfe01;
			16'head9: y = 16'hfe01;
			16'heada: y = 16'hfe01;
			16'headb: y = 16'hfe01;
			16'headc: y = 16'hfe01;
			16'headd: y = 16'hfe01;
			16'heade: y = 16'hfe01;
			16'headf: y = 16'hfe01;
			16'heae0: y = 16'hfe01;
			16'heae1: y = 16'hfe01;
			16'heae2: y = 16'hfe01;
			16'heae3: y = 16'hfe01;
			16'heae4: y = 16'hfe01;
			16'heae5: y = 16'hfe01;
			16'heae6: y = 16'hfe01;
			16'heae7: y = 16'hfe01;
			16'heae8: y = 16'hfe01;
			16'heae9: y = 16'hfe01;
			16'heaea: y = 16'hfe01;
			16'heaeb: y = 16'hfe01;
			16'heaec: y = 16'hfe01;
			16'heaed: y = 16'hfe01;
			16'heaee: y = 16'hfe01;
			16'heaef: y = 16'hfe01;
			16'heaf0: y = 16'hfe01;
			16'heaf1: y = 16'hfe01;
			16'heaf2: y = 16'hfe01;
			16'heaf3: y = 16'hfe01;
			16'heaf4: y = 16'hfe01;
			16'heaf5: y = 16'hfe01;
			16'heaf6: y = 16'hfe01;
			16'heaf7: y = 16'hfe01;
			16'heaf8: y = 16'hfe01;
			16'heaf9: y = 16'hfe01;
			16'heafa: y = 16'hfe01;
			16'heafb: y = 16'hfe01;
			16'heafc: y = 16'hfe01;
			16'heafd: y = 16'hfe01;
			16'heafe: y = 16'hfe01;
			16'heaff: y = 16'hfe01;
			16'heb00: y = 16'hfe01;
			16'heb01: y = 16'hfe01;
			16'heb02: y = 16'hfe01;
			16'heb03: y = 16'hfe01;
			16'heb04: y = 16'hfe01;
			16'heb05: y = 16'hfe01;
			16'heb06: y = 16'hfe01;
			16'heb07: y = 16'hfe01;
			16'heb08: y = 16'hfe01;
			16'heb09: y = 16'hfe01;
			16'heb0a: y = 16'hfe01;
			16'heb0b: y = 16'hfe01;
			16'heb0c: y = 16'hfe01;
			16'heb0d: y = 16'hfe01;
			16'heb0e: y = 16'hfe01;
			16'heb0f: y = 16'hfe01;
			16'heb10: y = 16'hfe01;
			16'heb11: y = 16'hfe01;
			16'heb12: y = 16'hfe01;
			16'heb13: y = 16'hfe01;
			16'heb14: y = 16'hfe01;
			16'heb15: y = 16'hfe01;
			16'heb16: y = 16'hfe01;
			16'heb17: y = 16'hfe01;
			16'heb18: y = 16'hfe01;
			16'heb19: y = 16'hfe01;
			16'heb1a: y = 16'hfe01;
			16'heb1b: y = 16'hfe01;
			16'heb1c: y = 16'hfe01;
			16'heb1d: y = 16'hfe01;
			16'heb1e: y = 16'hfe01;
			16'heb1f: y = 16'hfe01;
			16'heb20: y = 16'hfe01;
			16'heb21: y = 16'hfe01;
			16'heb22: y = 16'hfe01;
			16'heb23: y = 16'hfe01;
			16'heb24: y = 16'hfe01;
			16'heb25: y = 16'hfe01;
			16'heb26: y = 16'hfe01;
			16'heb27: y = 16'hfe01;
			16'heb28: y = 16'hfe01;
			16'heb29: y = 16'hfe01;
			16'heb2a: y = 16'hfe01;
			16'heb2b: y = 16'hfe01;
			16'heb2c: y = 16'hfe01;
			16'heb2d: y = 16'hfe01;
			16'heb2e: y = 16'hfe01;
			16'heb2f: y = 16'hfe01;
			16'heb30: y = 16'hfe01;
			16'heb31: y = 16'hfe01;
			16'heb32: y = 16'hfe01;
			16'heb33: y = 16'hfe01;
			16'heb34: y = 16'hfe01;
			16'heb35: y = 16'hfe01;
			16'heb36: y = 16'hfe01;
			16'heb37: y = 16'hfe01;
			16'heb38: y = 16'hfe01;
			16'heb39: y = 16'hfe01;
			16'heb3a: y = 16'hfe01;
			16'heb3b: y = 16'hfe01;
			16'heb3c: y = 16'hfe01;
			16'heb3d: y = 16'hfe01;
			16'heb3e: y = 16'hfe01;
			16'heb3f: y = 16'hfe01;
			16'heb40: y = 16'hfe01;
			16'heb41: y = 16'hfe01;
			16'heb42: y = 16'hfe01;
			16'heb43: y = 16'hfe01;
			16'heb44: y = 16'hfe01;
			16'heb45: y = 16'hfe01;
			16'heb46: y = 16'hfe01;
			16'heb47: y = 16'hfe01;
			16'heb48: y = 16'hfe01;
			16'heb49: y = 16'hfe01;
			16'heb4a: y = 16'hfe01;
			16'heb4b: y = 16'hfe01;
			16'heb4c: y = 16'hfe01;
			16'heb4d: y = 16'hfe01;
			16'heb4e: y = 16'hfe01;
			16'heb4f: y = 16'hfe01;
			16'heb50: y = 16'hfe01;
			16'heb51: y = 16'hfe01;
			16'heb52: y = 16'hfe01;
			16'heb53: y = 16'hfe01;
			16'heb54: y = 16'hfe01;
			16'heb55: y = 16'hfe01;
			16'heb56: y = 16'hfe01;
			16'heb57: y = 16'hfe01;
			16'heb58: y = 16'hfe01;
			16'heb59: y = 16'hfe01;
			16'heb5a: y = 16'hfe01;
			16'heb5b: y = 16'hfe01;
			16'heb5c: y = 16'hfe01;
			16'heb5d: y = 16'hfe01;
			16'heb5e: y = 16'hfe01;
			16'heb5f: y = 16'hfe01;
			16'heb60: y = 16'hfe01;
			16'heb61: y = 16'hfe01;
			16'heb62: y = 16'hfe01;
			16'heb63: y = 16'hfe01;
			16'heb64: y = 16'hfe01;
			16'heb65: y = 16'hfe01;
			16'heb66: y = 16'hfe01;
			16'heb67: y = 16'hfe01;
			16'heb68: y = 16'hfe01;
			16'heb69: y = 16'hfe01;
			16'heb6a: y = 16'hfe01;
			16'heb6b: y = 16'hfe01;
			16'heb6c: y = 16'hfe01;
			16'heb6d: y = 16'hfe01;
			16'heb6e: y = 16'hfe01;
			16'heb6f: y = 16'hfe01;
			16'heb70: y = 16'hfe01;
			16'heb71: y = 16'hfe01;
			16'heb72: y = 16'hfe01;
			16'heb73: y = 16'hfe01;
			16'heb74: y = 16'hfe01;
			16'heb75: y = 16'hfe01;
			16'heb76: y = 16'hfe01;
			16'heb77: y = 16'hfe01;
			16'heb78: y = 16'hfe01;
			16'heb79: y = 16'hfe01;
			16'heb7a: y = 16'hfe01;
			16'heb7b: y = 16'hfe01;
			16'heb7c: y = 16'hfe01;
			16'heb7d: y = 16'hfe01;
			16'heb7e: y = 16'hfe01;
			16'heb7f: y = 16'hfe01;
			16'heb80: y = 16'hfe01;
			16'heb81: y = 16'hfe01;
			16'heb82: y = 16'hfe01;
			16'heb83: y = 16'hfe01;
			16'heb84: y = 16'hfe01;
			16'heb85: y = 16'hfe01;
			16'heb86: y = 16'hfe01;
			16'heb87: y = 16'hfe01;
			16'heb88: y = 16'hfe01;
			16'heb89: y = 16'hfe01;
			16'heb8a: y = 16'hfe01;
			16'heb8b: y = 16'hfe01;
			16'heb8c: y = 16'hfe01;
			16'heb8d: y = 16'hfe01;
			16'heb8e: y = 16'hfe01;
			16'heb8f: y = 16'hfe01;
			16'heb90: y = 16'hfe01;
			16'heb91: y = 16'hfe01;
			16'heb92: y = 16'hfe01;
			16'heb93: y = 16'hfe01;
			16'heb94: y = 16'hfe01;
			16'heb95: y = 16'hfe01;
			16'heb96: y = 16'hfe01;
			16'heb97: y = 16'hfe01;
			16'heb98: y = 16'hfe01;
			16'heb99: y = 16'hfe01;
			16'heb9a: y = 16'hfe01;
			16'heb9b: y = 16'hfe01;
			16'heb9c: y = 16'hfe01;
			16'heb9d: y = 16'hfe01;
			16'heb9e: y = 16'hfe01;
			16'heb9f: y = 16'hfe01;
			16'heba0: y = 16'hfe01;
			16'heba1: y = 16'hfe01;
			16'heba2: y = 16'hfe01;
			16'heba3: y = 16'hfe01;
			16'heba4: y = 16'hfe01;
			16'heba5: y = 16'hfe01;
			16'heba6: y = 16'hfe01;
			16'heba7: y = 16'hfe01;
			16'heba8: y = 16'hfe01;
			16'heba9: y = 16'hfe01;
			16'hebaa: y = 16'hfe01;
			16'hebab: y = 16'hfe01;
			16'hebac: y = 16'hfe01;
			16'hebad: y = 16'hfe01;
			16'hebae: y = 16'hfe01;
			16'hebaf: y = 16'hfe01;
			16'hebb0: y = 16'hfe01;
			16'hebb1: y = 16'hfe01;
			16'hebb2: y = 16'hfe01;
			16'hebb3: y = 16'hfe01;
			16'hebb4: y = 16'hfe01;
			16'hebb5: y = 16'hfe01;
			16'hebb6: y = 16'hfe01;
			16'hebb7: y = 16'hfe01;
			16'hebb8: y = 16'hfe01;
			16'hebb9: y = 16'hfe01;
			16'hebba: y = 16'hfe01;
			16'hebbb: y = 16'hfe01;
			16'hebbc: y = 16'hfe01;
			16'hebbd: y = 16'hfe01;
			16'hebbe: y = 16'hfe01;
			16'hebbf: y = 16'hfe01;
			16'hebc0: y = 16'hfe01;
			16'hebc1: y = 16'hfe01;
			16'hebc2: y = 16'hfe01;
			16'hebc3: y = 16'hfe01;
			16'hebc4: y = 16'hfe01;
			16'hebc5: y = 16'hfe01;
			16'hebc6: y = 16'hfe01;
			16'hebc7: y = 16'hfe01;
			16'hebc8: y = 16'hfe01;
			16'hebc9: y = 16'hfe01;
			16'hebca: y = 16'hfe01;
			16'hebcb: y = 16'hfe01;
			16'hebcc: y = 16'hfe01;
			16'hebcd: y = 16'hfe01;
			16'hebce: y = 16'hfe01;
			16'hebcf: y = 16'hfe01;
			16'hebd0: y = 16'hfe01;
			16'hebd1: y = 16'hfe01;
			16'hebd2: y = 16'hfe01;
			16'hebd3: y = 16'hfe01;
			16'hebd4: y = 16'hfe01;
			16'hebd5: y = 16'hfe01;
			16'hebd6: y = 16'hfe01;
			16'hebd7: y = 16'hfe01;
			16'hebd8: y = 16'hfe01;
			16'hebd9: y = 16'hfe01;
			16'hebda: y = 16'hfe01;
			16'hebdb: y = 16'hfe01;
			16'hebdc: y = 16'hfe01;
			16'hebdd: y = 16'hfe01;
			16'hebde: y = 16'hfe01;
			16'hebdf: y = 16'hfe01;
			16'hebe0: y = 16'hfe01;
			16'hebe1: y = 16'hfe01;
			16'hebe2: y = 16'hfe01;
			16'hebe3: y = 16'hfe01;
			16'hebe4: y = 16'hfe01;
			16'hebe5: y = 16'hfe01;
			16'hebe6: y = 16'hfe01;
			16'hebe7: y = 16'hfe01;
			16'hebe8: y = 16'hfe01;
			16'hebe9: y = 16'hfe01;
			16'hebea: y = 16'hfe01;
			16'hebeb: y = 16'hfe01;
			16'hebec: y = 16'hfe01;
			16'hebed: y = 16'hfe01;
			16'hebee: y = 16'hfe01;
			16'hebef: y = 16'hfe01;
			16'hebf0: y = 16'hfe01;
			16'hebf1: y = 16'hfe01;
			16'hebf2: y = 16'hfe01;
			16'hebf3: y = 16'hfe01;
			16'hebf4: y = 16'hfe01;
			16'hebf5: y = 16'hfe01;
			16'hebf6: y = 16'hfe01;
			16'hebf7: y = 16'hfe01;
			16'hebf8: y = 16'hfe01;
			16'hebf9: y = 16'hfe01;
			16'hebfa: y = 16'hfe01;
			16'hebfb: y = 16'hfe01;
			16'hebfc: y = 16'hfe01;
			16'hebfd: y = 16'hfe01;
			16'hebfe: y = 16'hfe01;
			16'hebff: y = 16'hfe01;
			16'hec00: y = 16'hfe01;
			16'hec01: y = 16'hfe01;
			16'hec02: y = 16'hfe01;
			16'hec03: y = 16'hfe01;
			16'hec04: y = 16'hfe01;
			16'hec05: y = 16'hfe01;
			16'hec06: y = 16'hfe01;
			16'hec07: y = 16'hfe01;
			16'hec08: y = 16'hfe01;
			16'hec09: y = 16'hfe01;
			16'hec0a: y = 16'hfe01;
			16'hec0b: y = 16'hfe01;
			16'hec0c: y = 16'hfe01;
			16'hec0d: y = 16'hfe01;
			16'hec0e: y = 16'hfe01;
			16'hec0f: y = 16'hfe01;
			16'hec10: y = 16'hfe01;
			16'hec11: y = 16'hfe01;
			16'hec12: y = 16'hfe01;
			16'hec13: y = 16'hfe01;
			16'hec14: y = 16'hfe01;
			16'hec15: y = 16'hfe01;
			16'hec16: y = 16'hfe01;
			16'hec17: y = 16'hfe01;
			16'hec18: y = 16'hfe01;
			16'hec19: y = 16'hfe01;
			16'hec1a: y = 16'hfe01;
			16'hec1b: y = 16'hfe01;
			16'hec1c: y = 16'hfe01;
			16'hec1d: y = 16'hfe01;
			16'hec1e: y = 16'hfe01;
			16'hec1f: y = 16'hfe01;
			16'hec20: y = 16'hfe01;
			16'hec21: y = 16'hfe01;
			16'hec22: y = 16'hfe01;
			16'hec23: y = 16'hfe01;
			16'hec24: y = 16'hfe01;
			16'hec25: y = 16'hfe01;
			16'hec26: y = 16'hfe01;
			16'hec27: y = 16'hfe01;
			16'hec28: y = 16'hfe01;
			16'hec29: y = 16'hfe01;
			16'hec2a: y = 16'hfe01;
			16'hec2b: y = 16'hfe01;
			16'hec2c: y = 16'hfe01;
			16'hec2d: y = 16'hfe01;
			16'hec2e: y = 16'hfe01;
			16'hec2f: y = 16'hfe01;
			16'hec30: y = 16'hfe01;
			16'hec31: y = 16'hfe01;
			16'hec32: y = 16'hfe01;
			16'hec33: y = 16'hfe01;
			16'hec34: y = 16'hfe01;
			16'hec35: y = 16'hfe01;
			16'hec36: y = 16'hfe01;
			16'hec37: y = 16'hfe01;
			16'hec38: y = 16'hfe01;
			16'hec39: y = 16'hfe01;
			16'hec3a: y = 16'hfe01;
			16'hec3b: y = 16'hfe01;
			16'hec3c: y = 16'hfe01;
			16'hec3d: y = 16'hfe01;
			16'hec3e: y = 16'hfe01;
			16'hec3f: y = 16'hfe01;
			16'hec40: y = 16'hfe01;
			16'hec41: y = 16'hfe01;
			16'hec42: y = 16'hfe01;
			16'hec43: y = 16'hfe01;
			16'hec44: y = 16'hfe01;
			16'hec45: y = 16'hfe01;
			16'hec46: y = 16'hfe01;
			16'hec47: y = 16'hfe01;
			16'hec48: y = 16'hfe01;
			16'hec49: y = 16'hfe01;
			16'hec4a: y = 16'hfe01;
			16'hec4b: y = 16'hfe01;
			16'hec4c: y = 16'hfe01;
			16'hec4d: y = 16'hfe01;
			16'hec4e: y = 16'hfe01;
			16'hec4f: y = 16'hfe01;
			16'hec50: y = 16'hfe01;
			16'hec51: y = 16'hfe01;
			16'hec52: y = 16'hfe01;
			16'hec53: y = 16'hfe01;
			16'hec54: y = 16'hfe01;
			16'hec55: y = 16'hfe01;
			16'hec56: y = 16'hfe01;
			16'hec57: y = 16'hfe01;
			16'hec58: y = 16'hfe01;
			16'hec59: y = 16'hfe01;
			16'hec5a: y = 16'hfe01;
			16'hec5b: y = 16'hfe01;
			16'hec5c: y = 16'hfe01;
			16'hec5d: y = 16'hfe01;
			16'hec5e: y = 16'hfe01;
			16'hec5f: y = 16'hfe01;
			16'hec60: y = 16'hfe01;
			16'hec61: y = 16'hfe01;
			16'hec62: y = 16'hfe01;
			16'hec63: y = 16'hfe01;
			16'hec64: y = 16'hfe01;
			16'hec65: y = 16'hfe01;
			16'hec66: y = 16'hfe01;
			16'hec67: y = 16'hfe01;
			16'hec68: y = 16'hfe01;
			16'hec69: y = 16'hfe01;
			16'hec6a: y = 16'hfe01;
			16'hec6b: y = 16'hfe01;
			16'hec6c: y = 16'hfe01;
			16'hec6d: y = 16'hfe01;
			16'hec6e: y = 16'hfe01;
			16'hec6f: y = 16'hfe01;
			16'hec70: y = 16'hfe01;
			16'hec71: y = 16'hfe01;
			16'hec72: y = 16'hfe01;
			16'hec73: y = 16'hfe01;
			16'hec74: y = 16'hfe01;
			16'hec75: y = 16'hfe01;
			16'hec76: y = 16'hfe01;
			16'hec77: y = 16'hfe01;
			16'hec78: y = 16'hfe01;
			16'hec79: y = 16'hfe01;
			16'hec7a: y = 16'hfe01;
			16'hec7b: y = 16'hfe01;
			16'hec7c: y = 16'hfe01;
			16'hec7d: y = 16'hfe01;
			16'hec7e: y = 16'hfe01;
			16'hec7f: y = 16'hfe01;
			16'hec80: y = 16'hfe01;
			16'hec81: y = 16'hfe01;
			16'hec82: y = 16'hfe01;
			16'hec83: y = 16'hfe01;
			16'hec84: y = 16'hfe01;
			16'hec85: y = 16'hfe01;
			16'hec86: y = 16'hfe01;
			16'hec87: y = 16'hfe01;
			16'hec88: y = 16'hfe01;
			16'hec89: y = 16'hfe01;
			16'hec8a: y = 16'hfe01;
			16'hec8b: y = 16'hfe01;
			16'hec8c: y = 16'hfe01;
			16'hec8d: y = 16'hfe01;
			16'hec8e: y = 16'hfe01;
			16'hec8f: y = 16'hfe01;
			16'hec90: y = 16'hfe01;
			16'hec91: y = 16'hfe01;
			16'hec92: y = 16'hfe01;
			16'hec93: y = 16'hfe01;
			16'hec94: y = 16'hfe01;
			16'hec95: y = 16'hfe01;
			16'hec96: y = 16'hfe01;
			16'hec97: y = 16'hfe01;
			16'hec98: y = 16'hfe01;
			16'hec99: y = 16'hfe01;
			16'hec9a: y = 16'hfe01;
			16'hec9b: y = 16'hfe01;
			16'hec9c: y = 16'hfe01;
			16'hec9d: y = 16'hfe01;
			16'hec9e: y = 16'hfe01;
			16'hec9f: y = 16'hfe01;
			16'heca0: y = 16'hfe01;
			16'heca1: y = 16'hfe01;
			16'heca2: y = 16'hfe01;
			16'heca3: y = 16'hfe01;
			16'heca4: y = 16'hfe01;
			16'heca5: y = 16'hfe01;
			16'heca6: y = 16'hfe01;
			16'heca7: y = 16'hfe01;
			16'heca8: y = 16'hfe01;
			16'heca9: y = 16'hfe01;
			16'hecaa: y = 16'hfe01;
			16'hecab: y = 16'hfe01;
			16'hecac: y = 16'hfe01;
			16'hecad: y = 16'hfe01;
			16'hecae: y = 16'hfe01;
			16'hecaf: y = 16'hfe01;
			16'hecb0: y = 16'hfe01;
			16'hecb1: y = 16'hfe01;
			16'hecb2: y = 16'hfe01;
			16'hecb3: y = 16'hfe01;
			16'hecb4: y = 16'hfe01;
			16'hecb5: y = 16'hfe01;
			16'hecb6: y = 16'hfe01;
			16'hecb7: y = 16'hfe01;
			16'hecb8: y = 16'hfe01;
			16'hecb9: y = 16'hfe01;
			16'hecba: y = 16'hfe01;
			16'hecbb: y = 16'hfe01;
			16'hecbc: y = 16'hfe01;
			16'hecbd: y = 16'hfe01;
			16'hecbe: y = 16'hfe01;
			16'hecbf: y = 16'hfe01;
			16'hecc0: y = 16'hfe01;
			16'hecc1: y = 16'hfe01;
			16'hecc2: y = 16'hfe01;
			16'hecc3: y = 16'hfe01;
			16'hecc4: y = 16'hfe01;
			16'hecc5: y = 16'hfe01;
			16'hecc6: y = 16'hfe01;
			16'hecc7: y = 16'hfe01;
			16'hecc8: y = 16'hfe01;
			16'hecc9: y = 16'hfe01;
			16'hecca: y = 16'hfe01;
			16'heccb: y = 16'hfe01;
			16'heccc: y = 16'hfe01;
			16'heccd: y = 16'hfe01;
			16'hecce: y = 16'hfe01;
			16'heccf: y = 16'hfe01;
			16'hecd0: y = 16'hfe01;
			16'hecd1: y = 16'hfe01;
			16'hecd2: y = 16'hfe01;
			16'hecd3: y = 16'hfe01;
			16'hecd4: y = 16'hfe01;
			16'hecd5: y = 16'hfe01;
			16'hecd6: y = 16'hfe01;
			16'hecd7: y = 16'hfe01;
			16'hecd8: y = 16'hfe01;
			16'hecd9: y = 16'hfe01;
			16'hecda: y = 16'hfe01;
			16'hecdb: y = 16'hfe01;
			16'hecdc: y = 16'hfe01;
			16'hecdd: y = 16'hfe01;
			16'hecde: y = 16'hfe01;
			16'hecdf: y = 16'hfe01;
			16'hece0: y = 16'hfe01;
			16'hece1: y = 16'hfe01;
			16'hece2: y = 16'hfe01;
			16'hece3: y = 16'hfe01;
			16'hece4: y = 16'hfe01;
			16'hece5: y = 16'hfe01;
			16'hece6: y = 16'hfe01;
			16'hece7: y = 16'hfe01;
			16'hece8: y = 16'hfe01;
			16'hece9: y = 16'hfe01;
			16'hecea: y = 16'hfe01;
			16'heceb: y = 16'hfe01;
			16'hecec: y = 16'hfe01;
			16'heced: y = 16'hfe01;
			16'hecee: y = 16'hfe01;
			16'hecef: y = 16'hfe01;
			16'hecf0: y = 16'hfe01;
			16'hecf1: y = 16'hfe01;
			16'hecf2: y = 16'hfe01;
			16'hecf3: y = 16'hfe01;
			16'hecf4: y = 16'hfe01;
			16'hecf5: y = 16'hfe01;
			16'hecf6: y = 16'hfe01;
			16'hecf7: y = 16'hfe01;
			16'hecf8: y = 16'hfe01;
			16'hecf9: y = 16'hfe01;
			16'hecfa: y = 16'hfe01;
			16'hecfb: y = 16'hfe01;
			16'hecfc: y = 16'hfe01;
			16'hecfd: y = 16'hfe01;
			16'hecfe: y = 16'hfe01;
			16'hecff: y = 16'hfe01;
			16'hed00: y = 16'hfe01;
			16'hed01: y = 16'hfe01;
			16'hed02: y = 16'hfe01;
			16'hed03: y = 16'hfe01;
			16'hed04: y = 16'hfe01;
			16'hed05: y = 16'hfe01;
			16'hed06: y = 16'hfe01;
			16'hed07: y = 16'hfe01;
			16'hed08: y = 16'hfe01;
			16'hed09: y = 16'hfe01;
			16'hed0a: y = 16'hfe01;
			16'hed0b: y = 16'hfe01;
			16'hed0c: y = 16'hfe01;
			16'hed0d: y = 16'hfe01;
			16'hed0e: y = 16'hfe01;
			16'hed0f: y = 16'hfe01;
			16'hed10: y = 16'hfe01;
			16'hed11: y = 16'hfe01;
			16'hed12: y = 16'hfe01;
			16'hed13: y = 16'hfe01;
			16'hed14: y = 16'hfe01;
			16'hed15: y = 16'hfe01;
			16'hed16: y = 16'hfe01;
			16'hed17: y = 16'hfe01;
			16'hed18: y = 16'hfe01;
			16'hed19: y = 16'hfe01;
			16'hed1a: y = 16'hfe01;
			16'hed1b: y = 16'hfe01;
			16'hed1c: y = 16'hfe01;
			16'hed1d: y = 16'hfe01;
			16'hed1e: y = 16'hfe01;
			16'hed1f: y = 16'hfe01;
			16'hed20: y = 16'hfe01;
			16'hed21: y = 16'hfe01;
			16'hed22: y = 16'hfe01;
			16'hed23: y = 16'hfe01;
			16'hed24: y = 16'hfe01;
			16'hed25: y = 16'hfe01;
			16'hed26: y = 16'hfe01;
			16'hed27: y = 16'hfe01;
			16'hed28: y = 16'hfe01;
			16'hed29: y = 16'hfe01;
			16'hed2a: y = 16'hfe01;
			16'hed2b: y = 16'hfe01;
			16'hed2c: y = 16'hfe01;
			16'hed2d: y = 16'hfe01;
			16'hed2e: y = 16'hfe01;
			16'hed2f: y = 16'hfe01;
			16'hed30: y = 16'hfe01;
			16'hed31: y = 16'hfe01;
			16'hed32: y = 16'hfe01;
			16'hed33: y = 16'hfe01;
			16'hed34: y = 16'hfe01;
			16'hed35: y = 16'hfe01;
			16'hed36: y = 16'hfe01;
			16'hed37: y = 16'hfe01;
			16'hed38: y = 16'hfe01;
			16'hed39: y = 16'hfe01;
			16'hed3a: y = 16'hfe01;
			16'hed3b: y = 16'hfe01;
			16'hed3c: y = 16'hfe01;
			16'hed3d: y = 16'hfe01;
			16'hed3e: y = 16'hfe01;
			16'hed3f: y = 16'hfe01;
			16'hed40: y = 16'hfe01;
			16'hed41: y = 16'hfe01;
			16'hed42: y = 16'hfe01;
			16'hed43: y = 16'hfe01;
			16'hed44: y = 16'hfe01;
			16'hed45: y = 16'hfe01;
			16'hed46: y = 16'hfe01;
			16'hed47: y = 16'hfe01;
			16'hed48: y = 16'hfe01;
			16'hed49: y = 16'hfe01;
			16'hed4a: y = 16'hfe01;
			16'hed4b: y = 16'hfe01;
			16'hed4c: y = 16'hfe01;
			16'hed4d: y = 16'hfe01;
			16'hed4e: y = 16'hfe01;
			16'hed4f: y = 16'hfe01;
			16'hed50: y = 16'hfe01;
			16'hed51: y = 16'hfe01;
			16'hed52: y = 16'hfe01;
			16'hed53: y = 16'hfe01;
			16'hed54: y = 16'hfe01;
			16'hed55: y = 16'hfe01;
			16'hed56: y = 16'hfe01;
			16'hed57: y = 16'hfe01;
			16'hed58: y = 16'hfe01;
			16'hed59: y = 16'hfe01;
			16'hed5a: y = 16'hfe01;
			16'hed5b: y = 16'hfe01;
			16'hed5c: y = 16'hfe01;
			16'hed5d: y = 16'hfe01;
			16'hed5e: y = 16'hfe01;
			16'hed5f: y = 16'hfe01;
			16'hed60: y = 16'hfe01;
			16'hed61: y = 16'hfe01;
			16'hed62: y = 16'hfe01;
			16'hed63: y = 16'hfe01;
			16'hed64: y = 16'hfe01;
			16'hed65: y = 16'hfe01;
			16'hed66: y = 16'hfe01;
			16'hed67: y = 16'hfe01;
			16'hed68: y = 16'hfe01;
			16'hed69: y = 16'hfe01;
			16'hed6a: y = 16'hfe01;
			16'hed6b: y = 16'hfe01;
			16'hed6c: y = 16'hfe01;
			16'hed6d: y = 16'hfe01;
			16'hed6e: y = 16'hfe01;
			16'hed6f: y = 16'hfe01;
			16'hed70: y = 16'hfe01;
			16'hed71: y = 16'hfe01;
			16'hed72: y = 16'hfe01;
			16'hed73: y = 16'hfe01;
			16'hed74: y = 16'hfe01;
			16'hed75: y = 16'hfe01;
			16'hed76: y = 16'hfe01;
			16'hed77: y = 16'hfe01;
			16'hed78: y = 16'hfe01;
			16'hed79: y = 16'hfe01;
			16'hed7a: y = 16'hfe01;
			16'hed7b: y = 16'hfe01;
			16'hed7c: y = 16'hfe01;
			16'hed7d: y = 16'hfe01;
			16'hed7e: y = 16'hfe01;
			16'hed7f: y = 16'hfe01;
			16'hed80: y = 16'hfe01;
			16'hed81: y = 16'hfe01;
			16'hed82: y = 16'hfe01;
			16'hed83: y = 16'hfe01;
			16'hed84: y = 16'hfe01;
			16'hed85: y = 16'hfe01;
			16'hed86: y = 16'hfe01;
			16'hed87: y = 16'hfe01;
			16'hed88: y = 16'hfe01;
			16'hed89: y = 16'hfe01;
			16'hed8a: y = 16'hfe01;
			16'hed8b: y = 16'hfe01;
			16'hed8c: y = 16'hfe01;
			16'hed8d: y = 16'hfe01;
			16'hed8e: y = 16'hfe01;
			16'hed8f: y = 16'hfe01;
			16'hed90: y = 16'hfe01;
			16'hed91: y = 16'hfe01;
			16'hed92: y = 16'hfe01;
			16'hed93: y = 16'hfe01;
			16'hed94: y = 16'hfe01;
			16'hed95: y = 16'hfe01;
			16'hed96: y = 16'hfe01;
			16'hed97: y = 16'hfe01;
			16'hed98: y = 16'hfe01;
			16'hed99: y = 16'hfe01;
			16'hed9a: y = 16'hfe01;
			16'hed9b: y = 16'hfe01;
			16'hed9c: y = 16'hfe01;
			16'hed9d: y = 16'hfe01;
			16'hed9e: y = 16'hfe01;
			16'hed9f: y = 16'hfe01;
			16'heda0: y = 16'hfe01;
			16'heda1: y = 16'hfe01;
			16'heda2: y = 16'hfe01;
			16'heda3: y = 16'hfe01;
			16'heda4: y = 16'hfe01;
			16'heda5: y = 16'hfe01;
			16'heda6: y = 16'hfe01;
			16'heda7: y = 16'hfe01;
			16'heda8: y = 16'hfe01;
			16'heda9: y = 16'hfe01;
			16'hedaa: y = 16'hfe01;
			16'hedab: y = 16'hfe01;
			16'hedac: y = 16'hfe01;
			16'hedad: y = 16'hfe01;
			16'hedae: y = 16'hfe01;
			16'hedaf: y = 16'hfe01;
			16'hedb0: y = 16'hfe01;
			16'hedb1: y = 16'hfe01;
			16'hedb2: y = 16'hfe01;
			16'hedb3: y = 16'hfe01;
			16'hedb4: y = 16'hfe01;
			16'hedb5: y = 16'hfe01;
			16'hedb6: y = 16'hfe01;
			16'hedb7: y = 16'hfe01;
			16'hedb8: y = 16'hfe01;
			16'hedb9: y = 16'hfe01;
			16'hedba: y = 16'hfe01;
			16'hedbb: y = 16'hfe01;
			16'hedbc: y = 16'hfe01;
			16'hedbd: y = 16'hfe01;
			16'hedbe: y = 16'hfe01;
			16'hedbf: y = 16'hfe01;
			16'hedc0: y = 16'hfe01;
			16'hedc1: y = 16'hfe01;
			16'hedc2: y = 16'hfe01;
			16'hedc3: y = 16'hfe01;
			16'hedc4: y = 16'hfe01;
			16'hedc5: y = 16'hfe01;
			16'hedc6: y = 16'hfe01;
			16'hedc7: y = 16'hfe01;
			16'hedc8: y = 16'hfe01;
			16'hedc9: y = 16'hfe01;
			16'hedca: y = 16'hfe01;
			16'hedcb: y = 16'hfe01;
			16'hedcc: y = 16'hfe01;
			16'hedcd: y = 16'hfe01;
			16'hedce: y = 16'hfe01;
			16'hedcf: y = 16'hfe01;
			16'hedd0: y = 16'hfe01;
			16'hedd1: y = 16'hfe01;
			16'hedd2: y = 16'hfe01;
			16'hedd3: y = 16'hfe01;
			16'hedd4: y = 16'hfe01;
			16'hedd5: y = 16'hfe01;
			16'hedd6: y = 16'hfe01;
			16'hedd7: y = 16'hfe01;
			16'hedd8: y = 16'hfe01;
			16'hedd9: y = 16'hfe01;
			16'hedda: y = 16'hfe01;
			16'heddb: y = 16'hfe01;
			16'heddc: y = 16'hfe01;
			16'heddd: y = 16'hfe01;
			16'hedde: y = 16'hfe01;
			16'heddf: y = 16'hfe01;
			16'hede0: y = 16'hfe01;
			16'hede1: y = 16'hfe01;
			16'hede2: y = 16'hfe01;
			16'hede3: y = 16'hfe01;
			16'hede4: y = 16'hfe01;
			16'hede5: y = 16'hfe01;
			16'hede6: y = 16'hfe01;
			16'hede7: y = 16'hfe01;
			16'hede8: y = 16'hfe01;
			16'hede9: y = 16'hfe01;
			16'hedea: y = 16'hfe01;
			16'hedeb: y = 16'hfe01;
			16'hedec: y = 16'hfe01;
			16'heded: y = 16'hfe01;
			16'hedee: y = 16'hfe01;
			16'hedef: y = 16'hfe01;
			16'hedf0: y = 16'hfe01;
			16'hedf1: y = 16'hfe01;
			16'hedf2: y = 16'hfe01;
			16'hedf3: y = 16'hfe01;
			16'hedf4: y = 16'hfe01;
			16'hedf5: y = 16'hfe01;
			16'hedf6: y = 16'hfe01;
			16'hedf7: y = 16'hfe01;
			16'hedf8: y = 16'hfe01;
			16'hedf9: y = 16'hfe01;
			16'hedfa: y = 16'hfe01;
			16'hedfb: y = 16'hfe01;
			16'hedfc: y = 16'hfe01;
			16'hedfd: y = 16'hfe01;
			16'hedfe: y = 16'hfe01;
			16'hedff: y = 16'hfe01;
			16'hee00: y = 16'hfe01;
			16'hee01: y = 16'hfe01;
			16'hee02: y = 16'hfe01;
			16'hee03: y = 16'hfe01;
			16'hee04: y = 16'hfe01;
			16'hee05: y = 16'hfe01;
			16'hee06: y = 16'hfe01;
			16'hee07: y = 16'hfe01;
			16'hee08: y = 16'hfe01;
			16'hee09: y = 16'hfe01;
			16'hee0a: y = 16'hfe01;
			16'hee0b: y = 16'hfe01;
			16'hee0c: y = 16'hfe01;
			16'hee0d: y = 16'hfe01;
			16'hee0e: y = 16'hfe01;
			16'hee0f: y = 16'hfe01;
			16'hee10: y = 16'hfe01;
			16'hee11: y = 16'hfe01;
			16'hee12: y = 16'hfe01;
			16'hee13: y = 16'hfe01;
			16'hee14: y = 16'hfe01;
			16'hee15: y = 16'hfe01;
			16'hee16: y = 16'hfe01;
			16'hee17: y = 16'hfe01;
			16'hee18: y = 16'hfe01;
			16'hee19: y = 16'hfe01;
			16'hee1a: y = 16'hfe01;
			16'hee1b: y = 16'hfe01;
			16'hee1c: y = 16'hfe01;
			16'hee1d: y = 16'hfe01;
			16'hee1e: y = 16'hfe01;
			16'hee1f: y = 16'hfe01;
			16'hee20: y = 16'hfe01;
			16'hee21: y = 16'hfe01;
			16'hee22: y = 16'hfe01;
			16'hee23: y = 16'hfe01;
			16'hee24: y = 16'hfe01;
			16'hee25: y = 16'hfe01;
			16'hee26: y = 16'hfe01;
			16'hee27: y = 16'hfe01;
			16'hee28: y = 16'hfe01;
			16'hee29: y = 16'hfe01;
			16'hee2a: y = 16'hfe01;
			16'hee2b: y = 16'hfe01;
			16'hee2c: y = 16'hfe01;
			16'hee2d: y = 16'hfe01;
			16'hee2e: y = 16'hfe01;
			16'hee2f: y = 16'hfe01;
			16'hee30: y = 16'hfe01;
			16'hee31: y = 16'hfe01;
			16'hee32: y = 16'hfe01;
			16'hee33: y = 16'hfe01;
			16'hee34: y = 16'hfe01;
			16'hee35: y = 16'hfe01;
			16'hee36: y = 16'hfe01;
			16'hee37: y = 16'hfe01;
			16'hee38: y = 16'hfe01;
			16'hee39: y = 16'hfe01;
			16'hee3a: y = 16'hfe01;
			16'hee3b: y = 16'hfe01;
			16'hee3c: y = 16'hfe01;
			16'hee3d: y = 16'hfe01;
			16'hee3e: y = 16'hfe01;
			16'hee3f: y = 16'hfe01;
			16'hee40: y = 16'hfe01;
			16'hee41: y = 16'hfe01;
			16'hee42: y = 16'hfe01;
			16'hee43: y = 16'hfe01;
			16'hee44: y = 16'hfe01;
			16'hee45: y = 16'hfe01;
			16'hee46: y = 16'hfe01;
			16'hee47: y = 16'hfe01;
			16'hee48: y = 16'hfe01;
			16'hee49: y = 16'hfe01;
			16'hee4a: y = 16'hfe01;
			16'hee4b: y = 16'hfe01;
			16'hee4c: y = 16'hfe01;
			16'hee4d: y = 16'hfe01;
			16'hee4e: y = 16'hfe01;
			16'hee4f: y = 16'hfe01;
			16'hee50: y = 16'hfe01;
			16'hee51: y = 16'hfe01;
			16'hee52: y = 16'hfe01;
			16'hee53: y = 16'hfe01;
			16'hee54: y = 16'hfe01;
			16'hee55: y = 16'hfe01;
			16'hee56: y = 16'hfe01;
			16'hee57: y = 16'hfe01;
			16'hee58: y = 16'hfe01;
			16'hee59: y = 16'hfe01;
			16'hee5a: y = 16'hfe01;
			16'hee5b: y = 16'hfe01;
			16'hee5c: y = 16'hfe01;
			16'hee5d: y = 16'hfe01;
			16'hee5e: y = 16'hfe01;
			16'hee5f: y = 16'hfe01;
			16'hee60: y = 16'hfe01;
			16'hee61: y = 16'hfe01;
			16'hee62: y = 16'hfe01;
			16'hee63: y = 16'hfe01;
			16'hee64: y = 16'hfe01;
			16'hee65: y = 16'hfe01;
			16'hee66: y = 16'hfe01;
			16'hee67: y = 16'hfe01;
			16'hee68: y = 16'hfe01;
			16'hee69: y = 16'hfe01;
			16'hee6a: y = 16'hfe01;
			16'hee6b: y = 16'hfe01;
			16'hee6c: y = 16'hfe01;
			16'hee6d: y = 16'hfe01;
			16'hee6e: y = 16'hfe01;
			16'hee6f: y = 16'hfe01;
			16'hee70: y = 16'hfe01;
			16'hee71: y = 16'hfe01;
			16'hee72: y = 16'hfe01;
			16'hee73: y = 16'hfe01;
			16'hee74: y = 16'hfe01;
			16'hee75: y = 16'hfe01;
			16'hee76: y = 16'hfe01;
			16'hee77: y = 16'hfe01;
			16'hee78: y = 16'hfe01;
			16'hee79: y = 16'hfe01;
			16'hee7a: y = 16'hfe01;
			16'hee7b: y = 16'hfe01;
			16'hee7c: y = 16'hfe01;
			16'hee7d: y = 16'hfe01;
			16'hee7e: y = 16'hfe01;
			16'hee7f: y = 16'hfe01;
			16'hee80: y = 16'hfe01;
			16'hee81: y = 16'hfe01;
			16'hee82: y = 16'hfe01;
			16'hee83: y = 16'hfe01;
			16'hee84: y = 16'hfe01;
			16'hee85: y = 16'hfe01;
			16'hee86: y = 16'hfe01;
			16'hee87: y = 16'hfe01;
			16'hee88: y = 16'hfe01;
			16'hee89: y = 16'hfe01;
			16'hee8a: y = 16'hfe01;
			16'hee8b: y = 16'hfe01;
			16'hee8c: y = 16'hfe01;
			16'hee8d: y = 16'hfe01;
			16'hee8e: y = 16'hfe01;
			16'hee8f: y = 16'hfe01;
			16'hee90: y = 16'hfe01;
			16'hee91: y = 16'hfe01;
			16'hee92: y = 16'hfe01;
			16'hee93: y = 16'hfe01;
			16'hee94: y = 16'hfe01;
			16'hee95: y = 16'hfe01;
			16'hee96: y = 16'hfe01;
			16'hee97: y = 16'hfe01;
			16'hee98: y = 16'hfe01;
			16'hee99: y = 16'hfe01;
			16'hee9a: y = 16'hfe01;
			16'hee9b: y = 16'hfe01;
			16'hee9c: y = 16'hfe01;
			16'hee9d: y = 16'hfe01;
			16'hee9e: y = 16'hfe01;
			16'hee9f: y = 16'hfe01;
			16'heea0: y = 16'hfe01;
			16'heea1: y = 16'hfe01;
			16'heea2: y = 16'hfe01;
			16'heea3: y = 16'hfe01;
			16'heea4: y = 16'hfe01;
			16'heea5: y = 16'hfe01;
			16'heea6: y = 16'hfe01;
			16'heea7: y = 16'hfe01;
			16'heea8: y = 16'hfe01;
			16'heea9: y = 16'hfe01;
			16'heeaa: y = 16'hfe01;
			16'heeab: y = 16'hfe01;
			16'heeac: y = 16'hfe01;
			16'heead: y = 16'hfe01;
			16'heeae: y = 16'hfe01;
			16'heeaf: y = 16'hfe01;
			16'heeb0: y = 16'hfe01;
			16'heeb1: y = 16'hfe01;
			16'heeb2: y = 16'hfe01;
			16'heeb3: y = 16'hfe01;
			16'heeb4: y = 16'hfe01;
			16'heeb5: y = 16'hfe01;
			16'heeb6: y = 16'hfe01;
			16'heeb7: y = 16'hfe01;
			16'heeb8: y = 16'hfe01;
			16'heeb9: y = 16'hfe01;
			16'heeba: y = 16'hfe01;
			16'heebb: y = 16'hfe01;
			16'heebc: y = 16'hfe01;
			16'heebd: y = 16'hfe01;
			16'heebe: y = 16'hfe01;
			16'heebf: y = 16'hfe01;
			16'heec0: y = 16'hfe01;
			16'heec1: y = 16'hfe01;
			16'heec2: y = 16'hfe01;
			16'heec3: y = 16'hfe01;
			16'heec4: y = 16'hfe01;
			16'heec5: y = 16'hfe01;
			16'heec6: y = 16'hfe01;
			16'heec7: y = 16'hfe01;
			16'heec8: y = 16'hfe01;
			16'heec9: y = 16'hfe01;
			16'heeca: y = 16'hfe01;
			16'heecb: y = 16'hfe01;
			16'heecc: y = 16'hfe01;
			16'heecd: y = 16'hfe01;
			16'heece: y = 16'hfe01;
			16'heecf: y = 16'hfe01;
			16'heed0: y = 16'hfe01;
			16'heed1: y = 16'hfe01;
			16'heed2: y = 16'hfe01;
			16'heed3: y = 16'hfe01;
			16'heed4: y = 16'hfe01;
			16'heed5: y = 16'hfe01;
			16'heed6: y = 16'hfe01;
			16'heed7: y = 16'hfe01;
			16'heed8: y = 16'hfe01;
			16'heed9: y = 16'hfe01;
			16'heeda: y = 16'hfe01;
			16'heedb: y = 16'hfe01;
			16'heedc: y = 16'hfe01;
			16'heedd: y = 16'hfe01;
			16'heede: y = 16'hfe01;
			16'heedf: y = 16'hfe01;
			16'heee0: y = 16'hfe01;
			16'heee1: y = 16'hfe01;
			16'heee2: y = 16'hfe01;
			16'heee3: y = 16'hfe01;
			16'heee4: y = 16'hfe01;
			16'heee5: y = 16'hfe01;
			16'heee6: y = 16'hfe01;
			16'heee7: y = 16'hfe01;
			16'heee8: y = 16'hfe01;
			16'heee9: y = 16'hfe01;
			16'heeea: y = 16'hfe01;
			16'heeeb: y = 16'hfe01;
			16'heeec: y = 16'hfe01;
			16'heeed: y = 16'hfe01;
			16'heeee: y = 16'hfe01;
			16'heeef: y = 16'hfe01;
			16'heef0: y = 16'hfe01;
			16'heef1: y = 16'hfe01;
			16'heef2: y = 16'hfe01;
			16'heef3: y = 16'hfe01;
			16'heef4: y = 16'hfe01;
			16'heef5: y = 16'hfe01;
			16'heef6: y = 16'hfe01;
			16'heef7: y = 16'hfe01;
			16'heef8: y = 16'hfe01;
			16'heef9: y = 16'hfe01;
			16'heefa: y = 16'hfe01;
			16'heefb: y = 16'hfe01;
			16'heefc: y = 16'hfe01;
			16'heefd: y = 16'hfe01;
			16'heefe: y = 16'hfe01;
			16'heeff: y = 16'hfe01;
			16'hef00: y = 16'hfe01;
			16'hef01: y = 16'hfe01;
			16'hef02: y = 16'hfe01;
			16'hef03: y = 16'hfe01;
			16'hef04: y = 16'hfe01;
			16'hef05: y = 16'hfe01;
			16'hef06: y = 16'hfe01;
			16'hef07: y = 16'hfe01;
			16'hef08: y = 16'hfe01;
			16'hef09: y = 16'hfe01;
			16'hef0a: y = 16'hfe01;
			16'hef0b: y = 16'hfe01;
			16'hef0c: y = 16'hfe01;
			16'hef0d: y = 16'hfe01;
			16'hef0e: y = 16'hfe01;
			16'hef0f: y = 16'hfe01;
			16'hef10: y = 16'hfe01;
			16'hef11: y = 16'hfe01;
			16'hef12: y = 16'hfe01;
			16'hef13: y = 16'hfe01;
			16'hef14: y = 16'hfe01;
			16'hef15: y = 16'hfe01;
			16'hef16: y = 16'hfe01;
			16'hef17: y = 16'hfe01;
			16'hef18: y = 16'hfe01;
			16'hef19: y = 16'hfe01;
			16'hef1a: y = 16'hfe01;
			16'hef1b: y = 16'hfe01;
			16'hef1c: y = 16'hfe01;
			16'hef1d: y = 16'hfe01;
			16'hef1e: y = 16'hfe01;
			16'hef1f: y = 16'hfe01;
			16'hef20: y = 16'hfe01;
			16'hef21: y = 16'hfe01;
			16'hef22: y = 16'hfe01;
			16'hef23: y = 16'hfe01;
			16'hef24: y = 16'hfe01;
			16'hef25: y = 16'hfe01;
			16'hef26: y = 16'hfe01;
			16'hef27: y = 16'hfe01;
			16'hef28: y = 16'hfe01;
			16'hef29: y = 16'hfe01;
			16'hef2a: y = 16'hfe01;
			16'hef2b: y = 16'hfe01;
			16'hef2c: y = 16'hfe01;
			16'hef2d: y = 16'hfe01;
			16'hef2e: y = 16'hfe01;
			16'hef2f: y = 16'hfe01;
			16'hef30: y = 16'hfe01;
			16'hef31: y = 16'hfe01;
			16'hef32: y = 16'hfe01;
			16'hef33: y = 16'hfe01;
			16'hef34: y = 16'hfe01;
			16'hef35: y = 16'hfe01;
			16'hef36: y = 16'hfe01;
			16'hef37: y = 16'hfe01;
			16'hef38: y = 16'hfe01;
			16'hef39: y = 16'hfe01;
			16'hef3a: y = 16'hfe01;
			16'hef3b: y = 16'hfe01;
			16'hef3c: y = 16'hfe01;
			16'hef3d: y = 16'hfe01;
			16'hef3e: y = 16'hfe01;
			16'hef3f: y = 16'hfe01;
			16'hef40: y = 16'hfe01;
			16'hef41: y = 16'hfe01;
			16'hef42: y = 16'hfe01;
			16'hef43: y = 16'hfe01;
			16'hef44: y = 16'hfe01;
			16'hef45: y = 16'hfe01;
			16'hef46: y = 16'hfe01;
			16'hef47: y = 16'hfe01;
			16'hef48: y = 16'hfe01;
			16'hef49: y = 16'hfe01;
			16'hef4a: y = 16'hfe01;
			16'hef4b: y = 16'hfe01;
			16'hef4c: y = 16'hfe01;
			16'hef4d: y = 16'hfe01;
			16'hef4e: y = 16'hfe01;
			16'hef4f: y = 16'hfe01;
			16'hef50: y = 16'hfe01;
			16'hef51: y = 16'hfe01;
			16'hef52: y = 16'hfe01;
			16'hef53: y = 16'hfe01;
			16'hef54: y = 16'hfe01;
			16'hef55: y = 16'hfe01;
			16'hef56: y = 16'hfe01;
			16'hef57: y = 16'hfe01;
			16'hef58: y = 16'hfe01;
			16'hef59: y = 16'hfe01;
			16'hef5a: y = 16'hfe01;
			16'hef5b: y = 16'hfe01;
			16'hef5c: y = 16'hfe01;
			16'hef5d: y = 16'hfe01;
			16'hef5e: y = 16'hfe01;
			16'hef5f: y = 16'hfe01;
			16'hef60: y = 16'hfe01;
			16'hef61: y = 16'hfe01;
			16'hef62: y = 16'hfe01;
			16'hef63: y = 16'hfe01;
			16'hef64: y = 16'hfe01;
			16'hef65: y = 16'hfe01;
			16'hef66: y = 16'hfe01;
			16'hef67: y = 16'hfe01;
			16'hef68: y = 16'hfe01;
			16'hef69: y = 16'hfe01;
			16'hef6a: y = 16'hfe01;
			16'hef6b: y = 16'hfe01;
			16'hef6c: y = 16'hfe01;
			16'hef6d: y = 16'hfe01;
			16'hef6e: y = 16'hfe01;
			16'hef6f: y = 16'hfe01;
			16'hef70: y = 16'hfe01;
			16'hef71: y = 16'hfe01;
			16'hef72: y = 16'hfe01;
			16'hef73: y = 16'hfe01;
			16'hef74: y = 16'hfe01;
			16'hef75: y = 16'hfe01;
			16'hef76: y = 16'hfe01;
			16'hef77: y = 16'hfe01;
			16'hef78: y = 16'hfe01;
			16'hef79: y = 16'hfe01;
			16'hef7a: y = 16'hfe01;
			16'hef7b: y = 16'hfe01;
			16'hef7c: y = 16'hfe01;
			16'hef7d: y = 16'hfe01;
			16'hef7e: y = 16'hfe01;
			16'hef7f: y = 16'hfe01;
			16'hef80: y = 16'hfe01;
			16'hef81: y = 16'hfe01;
			16'hef82: y = 16'hfe01;
			16'hef83: y = 16'hfe01;
			16'hef84: y = 16'hfe01;
			16'hef85: y = 16'hfe01;
			16'hef86: y = 16'hfe01;
			16'hef87: y = 16'hfe01;
			16'hef88: y = 16'hfe01;
			16'hef89: y = 16'hfe01;
			16'hef8a: y = 16'hfe01;
			16'hef8b: y = 16'hfe01;
			16'hef8c: y = 16'hfe01;
			16'hef8d: y = 16'hfe01;
			16'hef8e: y = 16'hfe01;
			16'hef8f: y = 16'hfe01;
			16'hef90: y = 16'hfe01;
			16'hef91: y = 16'hfe01;
			16'hef92: y = 16'hfe01;
			16'hef93: y = 16'hfe01;
			16'hef94: y = 16'hfe01;
			16'hef95: y = 16'hfe01;
			16'hef96: y = 16'hfe01;
			16'hef97: y = 16'hfe01;
			16'hef98: y = 16'hfe01;
			16'hef99: y = 16'hfe01;
			16'hef9a: y = 16'hfe01;
			16'hef9b: y = 16'hfe01;
			16'hef9c: y = 16'hfe01;
			16'hef9d: y = 16'hfe01;
			16'hef9e: y = 16'hfe01;
			16'hef9f: y = 16'hfe01;
			16'hefa0: y = 16'hfe01;
			16'hefa1: y = 16'hfe01;
			16'hefa2: y = 16'hfe01;
			16'hefa3: y = 16'hfe01;
			16'hefa4: y = 16'hfe01;
			16'hefa5: y = 16'hfe01;
			16'hefa6: y = 16'hfe01;
			16'hefa7: y = 16'hfe01;
			16'hefa8: y = 16'hfe01;
			16'hefa9: y = 16'hfe01;
			16'hefaa: y = 16'hfe01;
			16'hefab: y = 16'hfe01;
			16'hefac: y = 16'hfe01;
			16'hefad: y = 16'hfe01;
			16'hefae: y = 16'hfe01;
			16'hefaf: y = 16'hfe01;
			16'hefb0: y = 16'hfe01;
			16'hefb1: y = 16'hfe01;
			16'hefb2: y = 16'hfe01;
			16'hefb3: y = 16'hfe01;
			16'hefb4: y = 16'hfe01;
			16'hefb5: y = 16'hfe01;
			16'hefb6: y = 16'hfe01;
			16'hefb7: y = 16'hfe01;
			16'hefb8: y = 16'hfe01;
			16'hefb9: y = 16'hfe01;
			16'hefba: y = 16'hfe01;
			16'hefbb: y = 16'hfe01;
			16'hefbc: y = 16'hfe01;
			16'hefbd: y = 16'hfe01;
			16'hefbe: y = 16'hfe01;
			16'hefbf: y = 16'hfe01;
			16'hefc0: y = 16'hfe01;
			16'hefc1: y = 16'hfe01;
			16'hefc2: y = 16'hfe01;
			16'hefc3: y = 16'hfe01;
			16'hefc4: y = 16'hfe01;
			16'hefc5: y = 16'hfe01;
			16'hefc6: y = 16'hfe01;
			16'hefc7: y = 16'hfe01;
			16'hefc8: y = 16'hfe01;
			16'hefc9: y = 16'hfe01;
			16'hefca: y = 16'hfe01;
			16'hefcb: y = 16'hfe01;
			16'hefcc: y = 16'hfe01;
			16'hefcd: y = 16'hfe01;
			16'hefce: y = 16'hfe01;
			16'hefcf: y = 16'hfe01;
			16'hefd0: y = 16'hfe01;
			16'hefd1: y = 16'hfe01;
			16'hefd2: y = 16'hfe01;
			16'hefd3: y = 16'hfe01;
			16'hefd4: y = 16'hfe01;
			16'hefd5: y = 16'hfe01;
			16'hefd6: y = 16'hfe01;
			16'hefd7: y = 16'hfe01;
			16'hefd8: y = 16'hfe01;
			16'hefd9: y = 16'hfe01;
			16'hefda: y = 16'hfe01;
			16'hefdb: y = 16'hfe01;
			16'hefdc: y = 16'hfe01;
			16'hefdd: y = 16'hfe01;
			16'hefde: y = 16'hfe01;
			16'hefdf: y = 16'hfe01;
			16'hefe0: y = 16'hfe01;
			16'hefe1: y = 16'hfe01;
			16'hefe2: y = 16'hfe01;
			16'hefe3: y = 16'hfe01;
			16'hefe4: y = 16'hfe01;
			16'hefe5: y = 16'hfe01;
			16'hefe6: y = 16'hfe01;
			16'hefe7: y = 16'hfe01;
			16'hefe8: y = 16'hfe01;
			16'hefe9: y = 16'hfe01;
			16'hefea: y = 16'hfe01;
			16'hefeb: y = 16'hfe01;
			16'hefec: y = 16'hfe01;
			16'hefed: y = 16'hfe01;
			16'hefee: y = 16'hfe01;
			16'hefef: y = 16'hfe01;
			16'heff0: y = 16'hfe01;
			16'heff1: y = 16'hfe01;
			16'heff2: y = 16'hfe01;
			16'heff3: y = 16'hfe01;
			16'heff4: y = 16'hfe01;
			16'heff5: y = 16'hfe01;
			16'heff6: y = 16'hfe01;
			16'heff7: y = 16'hfe01;
			16'heff8: y = 16'hfe01;
			16'heff9: y = 16'hfe01;
			16'heffa: y = 16'hfe01;
			16'heffb: y = 16'hfe01;
			16'heffc: y = 16'hfe01;
			16'heffd: y = 16'hfe01;
			16'heffe: y = 16'hfe01;
			16'hefff: y = 16'hfe01;
			16'hf000: y = 16'hfe01;
			16'hf001: y = 16'hfe01;
			16'hf002: y = 16'hfe01;
			16'hf003: y = 16'hfe01;
			16'hf004: y = 16'hfe01;
			16'hf005: y = 16'hfe01;
			16'hf006: y = 16'hfe01;
			16'hf007: y = 16'hfe01;
			16'hf008: y = 16'hfe01;
			16'hf009: y = 16'hfe01;
			16'hf00a: y = 16'hfe01;
			16'hf00b: y = 16'hfe01;
			16'hf00c: y = 16'hfe01;
			16'hf00d: y = 16'hfe01;
			16'hf00e: y = 16'hfe01;
			16'hf00f: y = 16'hfe01;
			16'hf010: y = 16'hfe01;
			16'hf011: y = 16'hfe01;
			16'hf012: y = 16'hfe01;
			16'hf013: y = 16'hfe01;
			16'hf014: y = 16'hfe01;
			16'hf015: y = 16'hfe01;
			16'hf016: y = 16'hfe01;
			16'hf017: y = 16'hfe01;
			16'hf018: y = 16'hfe01;
			16'hf019: y = 16'hfe01;
			16'hf01a: y = 16'hfe01;
			16'hf01b: y = 16'hfe01;
			16'hf01c: y = 16'hfe01;
			16'hf01d: y = 16'hfe01;
			16'hf01e: y = 16'hfe01;
			16'hf01f: y = 16'hfe01;
			16'hf020: y = 16'hfe01;
			16'hf021: y = 16'hfe01;
			16'hf022: y = 16'hfe01;
			16'hf023: y = 16'hfe01;
			16'hf024: y = 16'hfe01;
			16'hf025: y = 16'hfe01;
			16'hf026: y = 16'hfe01;
			16'hf027: y = 16'hfe01;
			16'hf028: y = 16'hfe01;
			16'hf029: y = 16'hfe01;
			16'hf02a: y = 16'hfe01;
			16'hf02b: y = 16'hfe01;
			16'hf02c: y = 16'hfe01;
			16'hf02d: y = 16'hfe01;
			16'hf02e: y = 16'hfe01;
			16'hf02f: y = 16'hfe01;
			16'hf030: y = 16'hfe01;
			16'hf031: y = 16'hfe01;
			16'hf032: y = 16'hfe01;
			16'hf033: y = 16'hfe01;
			16'hf034: y = 16'hfe01;
			16'hf035: y = 16'hfe01;
			16'hf036: y = 16'hfe01;
			16'hf037: y = 16'hfe01;
			16'hf038: y = 16'hfe01;
			16'hf039: y = 16'hfe01;
			16'hf03a: y = 16'hfe01;
			16'hf03b: y = 16'hfe01;
			16'hf03c: y = 16'hfe01;
			16'hf03d: y = 16'hfe01;
			16'hf03e: y = 16'hfe01;
			16'hf03f: y = 16'hfe01;
			16'hf040: y = 16'hfe01;
			16'hf041: y = 16'hfe01;
			16'hf042: y = 16'hfe01;
			16'hf043: y = 16'hfe01;
			16'hf044: y = 16'hfe01;
			16'hf045: y = 16'hfe01;
			16'hf046: y = 16'hfe01;
			16'hf047: y = 16'hfe01;
			16'hf048: y = 16'hfe01;
			16'hf049: y = 16'hfe01;
			16'hf04a: y = 16'hfe01;
			16'hf04b: y = 16'hfe01;
			16'hf04c: y = 16'hfe01;
			16'hf04d: y = 16'hfe01;
			16'hf04e: y = 16'hfe01;
			16'hf04f: y = 16'hfe01;
			16'hf050: y = 16'hfe01;
			16'hf051: y = 16'hfe01;
			16'hf052: y = 16'hfe01;
			16'hf053: y = 16'hfe01;
			16'hf054: y = 16'hfe01;
			16'hf055: y = 16'hfe01;
			16'hf056: y = 16'hfe01;
			16'hf057: y = 16'hfe01;
			16'hf058: y = 16'hfe01;
			16'hf059: y = 16'hfe01;
			16'hf05a: y = 16'hfe01;
			16'hf05b: y = 16'hfe01;
			16'hf05c: y = 16'hfe01;
			16'hf05d: y = 16'hfe01;
			16'hf05e: y = 16'hfe01;
			16'hf05f: y = 16'hfe01;
			16'hf060: y = 16'hfe01;
			16'hf061: y = 16'hfe01;
			16'hf062: y = 16'hfe01;
			16'hf063: y = 16'hfe01;
			16'hf064: y = 16'hfe01;
			16'hf065: y = 16'hfe01;
			16'hf066: y = 16'hfe01;
			16'hf067: y = 16'hfe01;
			16'hf068: y = 16'hfe01;
			16'hf069: y = 16'hfe01;
			16'hf06a: y = 16'hfe01;
			16'hf06b: y = 16'hfe01;
			16'hf06c: y = 16'hfe01;
			16'hf06d: y = 16'hfe01;
			16'hf06e: y = 16'hfe01;
			16'hf06f: y = 16'hfe01;
			16'hf070: y = 16'hfe01;
			16'hf071: y = 16'hfe01;
			16'hf072: y = 16'hfe01;
			16'hf073: y = 16'hfe01;
			16'hf074: y = 16'hfe01;
			16'hf075: y = 16'hfe01;
			16'hf076: y = 16'hfe01;
			16'hf077: y = 16'hfe01;
			16'hf078: y = 16'hfe01;
			16'hf079: y = 16'hfe01;
			16'hf07a: y = 16'hfe01;
			16'hf07b: y = 16'hfe01;
			16'hf07c: y = 16'hfe01;
			16'hf07d: y = 16'hfe01;
			16'hf07e: y = 16'hfe01;
			16'hf07f: y = 16'hfe01;
			16'hf080: y = 16'hfe01;
			16'hf081: y = 16'hfe01;
			16'hf082: y = 16'hfe01;
			16'hf083: y = 16'hfe01;
			16'hf084: y = 16'hfe01;
			16'hf085: y = 16'hfe01;
			16'hf086: y = 16'hfe01;
			16'hf087: y = 16'hfe01;
			16'hf088: y = 16'hfe01;
			16'hf089: y = 16'hfe01;
			16'hf08a: y = 16'hfe01;
			16'hf08b: y = 16'hfe01;
			16'hf08c: y = 16'hfe01;
			16'hf08d: y = 16'hfe01;
			16'hf08e: y = 16'hfe01;
			16'hf08f: y = 16'hfe01;
			16'hf090: y = 16'hfe01;
			16'hf091: y = 16'hfe01;
			16'hf092: y = 16'hfe01;
			16'hf093: y = 16'hfe01;
			16'hf094: y = 16'hfe01;
			16'hf095: y = 16'hfe01;
			16'hf096: y = 16'hfe01;
			16'hf097: y = 16'hfe01;
			16'hf098: y = 16'hfe01;
			16'hf099: y = 16'hfe01;
			16'hf09a: y = 16'hfe01;
			16'hf09b: y = 16'hfe01;
			16'hf09c: y = 16'hfe01;
			16'hf09d: y = 16'hfe01;
			16'hf09e: y = 16'hfe01;
			16'hf09f: y = 16'hfe01;
			16'hf0a0: y = 16'hfe01;
			16'hf0a1: y = 16'hfe01;
			16'hf0a2: y = 16'hfe01;
			16'hf0a3: y = 16'hfe01;
			16'hf0a4: y = 16'hfe01;
			16'hf0a5: y = 16'hfe01;
			16'hf0a6: y = 16'hfe01;
			16'hf0a7: y = 16'hfe01;
			16'hf0a8: y = 16'hfe01;
			16'hf0a9: y = 16'hfe01;
			16'hf0aa: y = 16'hfe01;
			16'hf0ab: y = 16'hfe01;
			16'hf0ac: y = 16'hfe01;
			16'hf0ad: y = 16'hfe01;
			16'hf0ae: y = 16'hfe01;
			16'hf0af: y = 16'hfe01;
			16'hf0b0: y = 16'hfe01;
			16'hf0b1: y = 16'hfe01;
			16'hf0b2: y = 16'hfe01;
			16'hf0b3: y = 16'hfe01;
			16'hf0b4: y = 16'hfe01;
			16'hf0b5: y = 16'hfe01;
			16'hf0b6: y = 16'hfe01;
			16'hf0b7: y = 16'hfe01;
			16'hf0b8: y = 16'hfe01;
			16'hf0b9: y = 16'hfe01;
			16'hf0ba: y = 16'hfe01;
			16'hf0bb: y = 16'hfe01;
			16'hf0bc: y = 16'hfe01;
			16'hf0bd: y = 16'hfe01;
			16'hf0be: y = 16'hfe01;
			16'hf0bf: y = 16'hfe01;
			16'hf0c0: y = 16'hfe01;
			16'hf0c1: y = 16'hfe01;
			16'hf0c2: y = 16'hfe01;
			16'hf0c3: y = 16'hfe01;
			16'hf0c4: y = 16'hfe01;
			16'hf0c5: y = 16'hfe01;
			16'hf0c6: y = 16'hfe01;
			16'hf0c7: y = 16'hfe01;
			16'hf0c8: y = 16'hfe01;
			16'hf0c9: y = 16'hfe01;
			16'hf0ca: y = 16'hfe01;
			16'hf0cb: y = 16'hfe01;
			16'hf0cc: y = 16'hfe01;
			16'hf0cd: y = 16'hfe01;
			16'hf0ce: y = 16'hfe01;
			16'hf0cf: y = 16'hfe01;
			16'hf0d0: y = 16'hfe01;
			16'hf0d1: y = 16'hfe01;
			16'hf0d2: y = 16'hfe01;
			16'hf0d3: y = 16'hfe01;
			16'hf0d4: y = 16'hfe01;
			16'hf0d5: y = 16'hfe01;
			16'hf0d6: y = 16'hfe01;
			16'hf0d7: y = 16'hfe01;
			16'hf0d8: y = 16'hfe01;
			16'hf0d9: y = 16'hfe01;
			16'hf0da: y = 16'hfe01;
			16'hf0db: y = 16'hfe01;
			16'hf0dc: y = 16'hfe01;
			16'hf0dd: y = 16'hfe01;
			16'hf0de: y = 16'hfe01;
			16'hf0df: y = 16'hfe01;
			16'hf0e0: y = 16'hfe01;
			16'hf0e1: y = 16'hfe01;
			16'hf0e2: y = 16'hfe01;
			16'hf0e3: y = 16'hfe01;
			16'hf0e4: y = 16'hfe01;
			16'hf0e5: y = 16'hfe01;
			16'hf0e6: y = 16'hfe01;
			16'hf0e7: y = 16'hfe01;
			16'hf0e8: y = 16'hfe01;
			16'hf0e9: y = 16'hfe01;
			16'hf0ea: y = 16'hfe01;
			16'hf0eb: y = 16'hfe01;
			16'hf0ec: y = 16'hfe01;
			16'hf0ed: y = 16'hfe01;
			16'hf0ee: y = 16'hfe01;
			16'hf0ef: y = 16'hfe01;
			16'hf0f0: y = 16'hfe01;
			16'hf0f1: y = 16'hfe01;
			16'hf0f2: y = 16'hfe01;
			16'hf0f3: y = 16'hfe01;
			16'hf0f4: y = 16'hfe01;
			16'hf0f5: y = 16'hfe01;
			16'hf0f6: y = 16'hfe01;
			16'hf0f7: y = 16'hfe01;
			16'hf0f8: y = 16'hfe01;
			16'hf0f9: y = 16'hfe01;
			16'hf0fa: y = 16'hfe01;
			16'hf0fb: y = 16'hfe01;
			16'hf0fc: y = 16'hfe01;
			16'hf0fd: y = 16'hfe01;
			16'hf0fe: y = 16'hfe01;
			16'hf0ff: y = 16'hfe01;
			16'hf100: y = 16'hfe01;
			16'hf101: y = 16'hfe01;
			16'hf102: y = 16'hfe01;
			16'hf103: y = 16'hfe01;
			16'hf104: y = 16'hfe01;
			16'hf105: y = 16'hfe01;
			16'hf106: y = 16'hfe01;
			16'hf107: y = 16'hfe01;
			16'hf108: y = 16'hfe01;
			16'hf109: y = 16'hfe01;
			16'hf10a: y = 16'hfe01;
			16'hf10b: y = 16'hfe01;
			16'hf10c: y = 16'hfe01;
			16'hf10d: y = 16'hfe01;
			16'hf10e: y = 16'hfe01;
			16'hf10f: y = 16'hfe01;
			16'hf110: y = 16'hfe01;
			16'hf111: y = 16'hfe01;
			16'hf112: y = 16'hfe01;
			16'hf113: y = 16'hfe01;
			16'hf114: y = 16'hfe01;
			16'hf115: y = 16'hfe01;
			16'hf116: y = 16'hfe01;
			16'hf117: y = 16'hfe01;
			16'hf118: y = 16'hfe01;
			16'hf119: y = 16'hfe01;
			16'hf11a: y = 16'hfe01;
			16'hf11b: y = 16'hfe01;
			16'hf11c: y = 16'hfe01;
			16'hf11d: y = 16'hfe01;
			16'hf11e: y = 16'hfe01;
			16'hf11f: y = 16'hfe01;
			16'hf120: y = 16'hfe01;
			16'hf121: y = 16'hfe01;
			16'hf122: y = 16'hfe01;
			16'hf123: y = 16'hfe01;
			16'hf124: y = 16'hfe01;
			16'hf125: y = 16'hfe01;
			16'hf126: y = 16'hfe01;
			16'hf127: y = 16'hfe01;
			16'hf128: y = 16'hfe01;
			16'hf129: y = 16'hfe01;
			16'hf12a: y = 16'hfe01;
			16'hf12b: y = 16'hfe01;
			16'hf12c: y = 16'hfe01;
			16'hf12d: y = 16'hfe01;
			16'hf12e: y = 16'hfe01;
			16'hf12f: y = 16'hfe01;
			16'hf130: y = 16'hfe01;
			16'hf131: y = 16'hfe01;
			16'hf132: y = 16'hfe01;
			16'hf133: y = 16'hfe01;
			16'hf134: y = 16'hfe01;
			16'hf135: y = 16'hfe01;
			16'hf136: y = 16'hfe01;
			16'hf137: y = 16'hfe01;
			16'hf138: y = 16'hfe01;
			16'hf139: y = 16'hfe01;
			16'hf13a: y = 16'hfe01;
			16'hf13b: y = 16'hfe01;
			16'hf13c: y = 16'hfe01;
			16'hf13d: y = 16'hfe01;
			16'hf13e: y = 16'hfe01;
			16'hf13f: y = 16'hfe01;
			16'hf140: y = 16'hfe01;
			16'hf141: y = 16'hfe01;
			16'hf142: y = 16'hfe01;
			16'hf143: y = 16'hfe01;
			16'hf144: y = 16'hfe01;
			16'hf145: y = 16'hfe01;
			16'hf146: y = 16'hfe01;
			16'hf147: y = 16'hfe01;
			16'hf148: y = 16'hfe01;
			16'hf149: y = 16'hfe01;
			16'hf14a: y = 16'hfe01;
			16'hf14b: y = 16'hfe01;
			16'hf14c: y = 16'hfe01;
			16'hf14d: y = 16'hfe01;
			16'hf14e: y = 16'hfe01;
			16'hf14f: y = 16'hfe01;
			16'hf150: y = 16'hfe01;
			16'hf151: y = 16'hfe01;
			16'hf152: y = 16'hfe01;
			16'hf153: y = 16'hfe01;
			16'hf154: y = 16'hfe01;
			16'hf155: y = 16'hfe01;
			16'hf156: y = 16'hfe01;
			16'hf157: y = 16'hfe01;
			16'hf158: y = 16'hfe01;
			16'hf159: y = 16'hfe01;
			16'hf15a: y = 16'hfe01;
			16'hf15b: y = 16'hfe01;
			16'hf15c: y = 16'hfe01;
			16'hf15d: y = 16'hfe01;
			16'hf15e: y = 16'hfe01;
			16'hf15f: y = 16'hfe01;
			16'hf160: y = 16'hfe01;
			16'hf161: y = 16'hfe01;
			16'hf162: y = 16'hfe01;
			16'hf163: y = 16'hfe01;
			16'hf164: y = 16'hfe01;
			16'hf165: y = 16'hfe01;
			16'hf166: y = 16'hfe01;
			16'hf167: y = 16'hfe01;
			16'hf168: y = 16'hfe01;
			16'hf169: y = 16'hfe01;
			16'hf16a: y = 16'hfe01;
			16'hf16b: y = 16'hfe01;
			16'hf16c: y = 16'hfe01;
			16'hf16d: y = 16'hfe01;
			16'hf16e: y = 16'hfe01;
			16'hf16f: y = 16'hfe01;
			16'hf170: y = 16'hfe01;
			16'hf171: y = 16'hfe01;
			16'hf172: y = 16'hfe01;
			16'hf173: y = 16'hfe01;
			16'hf174: y = 16'hfe01;
			16'hf175: y = 16'hfe01;
			16'hf176: y = 16'hfe01;
			16'hf177: y = 16'hfe01;
			16'hf178: y = 16'hfe01;
			16'hf179: y = 16'hfe01;
			16'hf17a: y = 16'hfe01;
			16'hf17b: y = 16'hfe01;
			16'hf17c: y = 16'hfe01;
			16'hf17d: y = 16'hfe01;
			16'hf17e: y = 16'hfe01;
			16'hf17f: y = 16'hfe01;
			16'hf180: y = 16'hfe01;
			16'hf181: y = 16'hfe01;
			16'hf182: y = 16'hfe01;
			16'hf183: y = 16'hfe01;
			16'hf184: y = 16'hfe01;
			16'hf185: y = 16'hfe01;
			16'hf186: y = 16'hfe01;
			16'hf187: y = 16'hfe01;
			16'hf188: y = 16'hfe01;
			16'hf189: y = 16'hfe01;
			16'hf18a: y = 16'hfe01;
			16'hf18b: y = 16'hfe01;
			16'hf18c: y = 16'hfe01;
			16'hf18d: y = 16'hfe01;
			16'hf18e: y = 16'hfe01;
			16'hf18f: y = 16'hfe01;
			16'hf190: y = 16'hfe01;
			16'hf191: y = 16'hfe01;
			16'hf192: y = 16'hfe01;
			16'hf193: y = 16'hfe01;
			16'hf194: y = 16'hfe01;
			16'hf195: y = 16'hfe01;
			16'hf196: y = 16'hfe01;
			16'hf197: y = 16'hfe01;
			16'hf198: y = 16'hfe01;
			16'hf199: y = 16'hfe01;
			16'hf19a: y = 16'hfe01;
			16'hf19b: y = 16'hfe01;
			16'hf19c: y = 16'hfe01;
			16'hf19d: y = 16'hfe01;
			16'hf19e: y = 16'hfe01;
			16'hf19f: y = 16'hfe01;
			16'hf1a0: y = 16'hfe01;
			16'hf1a1: y = 16'hfe01;
			16'hf1a2: y = 16'hfe01;
			16'hf1a3: y = 16'hfe01;
			16'hf1a4: y = 16'hfe01;
			16'hf1a5: y = 16'hfe01;
			16'hf1a6: y = 16'hfe01;
			16'hf1a7: y = 16'hfe01;
			16'hf1a8: y = 16'hfe01;
			16'hf1a9: y = 16'hfe01;
			16'hf1aa: y = 16'hfe01;
			16'hf1ab: y = 16'hfe01;
			16'hf1ac: y = 16'hfe01;
			16'hf1ad: y = 16'hfe01;
			16'hf1ae: y = 16'hfe01;
			16'hf1af: y = 16'hfe01;
			16'hf1b0: y = 16'hfe01;
			16'hf1b1: y = 16'hfe01;
			16'hf1b2: y = 16'hfe01;
			16'hf1b3: y = 16'hfe01;
			16'hf1b4: y = 16'hfe01;
			16'hf1b5: y = 16'hfe01;
			16'hf1b6: y = 16'hfe01;
			16'hf1b7: y = 16'hfe01;
			16'hf1b8: y = 16'hfe01;
			16'hf1b9: y = 16'hfe01;
			16'hf1ba: y = 16'hfe01;
			16'hf1bb: y = 16'hfe01;
			16'hf1bc: y = 16'hfe01;
			16'hf1bd: y = 16'hfe01;
			16'hf1be: y = 16'hfe01;
			16'hf1bf: y = 16'hfe01;
			16'hf1c0: y = 16'hfe01;
			16'hf1c1: y = 16'hfe01;
			16'hf1c2: y = 16'hfe01;
			16'hf1c3: y = 16'hfe01;
			16'hf1c4: y = 16'hfe01;
			16'hf1c5: y = 16'hfe01;
			16'hf1c6: y = 16'hfe01;
			16'hf1c7: y = 16'hfe01;
			16'hf1c8: y = 16'hfe01;
			16'hf1c9: y = 16'hfe01;
			16'hf1ca: y = 16'hfe01;
			16'hf1cb: y = 16'hfe01;
			16'hf1cc: y = 16'hfe01;
			16'hf1cd: y = 16'hfe01;
			16'hf1ce: y = 16'hfe01;
			16'hf1cf: y = 16'hfe01;
			16'hf1d0: y = 16'hfe01;
			16'hf1d1: y = 16'hfe01;
			16'hf1d2: y = 16'hfe01;
			16'hf1d3: y = 16'hfe01;
			16'hf1d4: y = 16'hfe01;
			16'hf1d5: y = 16'hfe01;
			16'hf1d6: y = 16'hfe01;
			16'hf1d7: y = 16'hfe01;
			16'hf1d8: y = 16'hfe01;
			16'hf1d9: y = 16'hfe01;
			16'hf1da: y = 16'hfe01;
			16'hf1db: y = 16'hfe01;
			16'hf1dc: y = 16'hfe01;
			16'hf1dd: y = 16'hfe01;
			16'hf1de: y = 16'hfe01;
			16'hf1df: y = 16'hfe01;
			16'hf1e0: y = 16'hfe01;
			16'hf1e1: y = 16'hfe01;
			16'hf1e2: y = 16'hfe01;
			16'hf1e3: y = 16'hfe01;
			16'hf1e4: y = 16'hfe01;
			16'hf1e5: y = 16'hfe01;
			16'hf1e6: y = 16'hfe01;
			16'hf1e7: y = 16'hfe01;
			16'hf1e8: y = 16'hfe01;
			16'hf1e9: y = 16'hfe01;
			16'hf1ea: y = 16'hfe01;
			16'hf1eb: y = 16'hfe01;
			16'hf1ec: y = 16'hfe01;
			16'hf1ed: y = 16'hfe01;
			16'hf1ee: y = 16'hfe01;
			16'hf1ef: y = 16'hfe01;
			16'hf1f0: y = 16'hfe01;
			16'hf1f1: y = 16'hfe01;
			16'hf1f2: y = 16'hfe01;
			16'hf1f3: y = 16'hfe01;
			16'hf1f4: y = 16'hfe01;
			16'hf1f5: y = 16'hfe01;
			16'hf1f6: y = 16'hfe01;
			16'hf1f7: y = 16'hfe01;
			16'hf1f8: y = 16'hfe01;
			16'hf1f9: y = 16'hfe01;
			16'hf1fa: y = 16'hfe01;
			16'hf1fb: y = 16'hfe01;
			16'hf1fc: y = 16'hfe01;
			16'hf1fd: y = 16'hfe01;
			16'hf1fe: y = 16'hfe01;
			16'hf1ff: y = 16'hfe01;
			16'hf200: y = 16'hfe01;
			16'hf201: y = 16'hfe01;
			16'hf202: y = 16'hfe01;
			16'hf203: y = 16'hfe01;
			16'hf204: y = 16'hfe01;
			16'hf205: y = 16'hfe01;
			16'hf206: y = 16'hfe01;
			16'hf207: y = 16'hfe01;
			16'hf208: y = 16'hfe01;
			16'hf209: y = 16'hfe01;
			16'hf20a: y = 16'hfe01;
			16'hf20b: y = 16'hfe01;
			16'hf20c: y = 16'hfe01;
			16'hf20d: y = 16'hfe01;
			16'hf20e: y = 16'hfe01;
			16'hf20f: y = 16'hfe01;
			16'hf210: y = 16'hfe01;
			16'hf211: y = 16'hfe01;
			16'hf212: y = 16'hfe01;
			16'hf213: y = 16'hfe01;
			16'hf214: y = 16'hfe01;
			16'hf215: y = 16'hfe01;
			16'hf216: y = 16'hfe01;
			16'hf217: y = 16'hfe01;
			16'hf218: y = 16'hfe01;
			16'hf219: y = 16'hfe01;
			16'hf21a: y = 16'hfe01;
			16'hf21b: y = 16'hfe01;
			16'hf21c: y = 16'hfe01;
			16'hf21d: y = 16'hfe01;
			16'hf21e: y = 16'hfe01;
			16'hf21f: y = 16'hfe01;
			16'hf220: y = 16'hfe01;
			16'hf221: y = 16'hfe01;
			16'hf222: y = 16'hfe01;
			16'hf223: y = 16'hfe01;
			16'hf224: y = 16'hfe01;
			16'hf225: y = 16'hfe01;
			16'hf226: y = 16'hfe01;
			16'hf227: y = 16'hfe01;
			16'hf228: y = 16'hfe01;
			16'hf229: y = 16'hfe01;
			16'hf22a: y = 16'hfe01;
			16'hf22b: y = 16'hfe01;
			16'hf22c: y = 16'hfe01;
			16'hf22d: y = 16'hfe01;
			16'hf22e: y = 16'hfe01;
			16'hf22f: y = 16'hfe01;
			16'hf230: y = 16'hfe01;
			16'hf231: y = 16'hfe01;
			16'hf232: y = 16'hfe01;
			16'hf233: y = 16'hfe01;
			16'hf234: y = 16'hfe01;
			16'hf235: y = 16'hfe01;
			16'hf236: y = 16'hfe01;
			16'hf237: y = 16'hfe01;
			16'hf238: y = 16'hfe01;
			16'hf239: y = 16'hfe01;
			16'hf23a: y = 16'hfe01;
			16'hf23b: y = 16'hfe01;
			16'hf23c: y = 16'hfe01;
			16'hf23d: y = 16'hfe01;
			16'hf23e: y = 16'hfe01;
			16'hf23f: y = 16'hfe01;
			16'hf240: y = 16'hfe01;
			16'hf241: y = 16'hfe01;
			16'hf242: y = 16'hfe01;
			16'hf243: y = 16'hfe01;
			16'hf244: y = 16'hfe01;
			16'hf245: y = 16'hfe01;
			16'hf246: y = 16'hfe01;
			16'hf247: y = 16'hfe01;
			16'hf248: y = 16'hfe01;
			16'hf249: y = 16'hfe01;
			16'hf24a: y = 16'hfe01;
			16'hf24b: y = 16'hfe01;
			16'hf24c: y = 16'hfe01;
			16'hf24d: y = 16'hfe01;
			16'hf24e: y = 16'hfe01;
			16'hf24f: y = 16'hfe01;
			16'hf250: y = 16'hfe01;
			16'hf251: y = 16'hfe01;
			16'hf252: y = 16'hfe01;
			16'hf253: y = 16'hfe01;
			16'hf254: y = 16'hfe01;
			16'hf255: y = 16'hfe01;
			16'hf256: y = 16'hfe01;
			16'hf257: y = 16'hfe01;
			16'hf258: y = 16'hfe01;
			16'hf259: y = 16'hfe01;
			16'hf25a: y = 16'hfe01;
			16'hf25b: y = 16'hfe01;
			16'hf25c: y = 16'hfe01;
			16'hf25d: y = 16'hfe01;
			16'hf25e: y = 16'hfe01;
			16'hf25f: y = 16'hfe01;
			16'hf260: y = 16'hfe01;
			16'hf261: y = 16'hfe01;
			16'hf262: y = 16'hfe01;
			16'hf263: y = 16'hfe01;
			16'hf264: y = 16'hfe01;
			16'hf265: y = 16'hfe01;
			16'hf266: y = 16'hfe01;
			16'hf267: y = 16'hfe01;
			16'hf268: y = 16'hfe01;
			16'hf269: y = 16'hfe01;
			16'hf26a: y = 16'hfe01;
			16'hf26b: y = 16'hfe01;
			16'hf26c: y = 16'hfe01;
			16'hf26d: y = 16'hfe01;
			16'hf26e: y = 16'hfe01;
			16'hf26f: y = 16'hfe01;
			16'hf270: y = 16'hfe01;
			16'hf271: y = 16'hfe01;
			16'hf272: y = 16'hfe01;
			16'hf273: y = 16'hfe01;
			16'hf274: y = 16'hfe01;
			16'hf275: y = 16'hfe01;
			16'hf276: y = 16'hfe01;
			16'hf277: y = 16'hfe01;
			16'hf278: y = 16'hfe01;
			16'hf279: y = 16'hfe01;
			16'hf27a: y = 16'hfe01;
			16'hf27b: y = 16'hfe01;
			16'hf27c: y = 16'hfe01;
			16'hf27d: y = 16'hfe01;
			16'hf27e: y = 16'hfe01;
			16'hf27f: y = 16'hfe01;
			16'hf280: y = 16'hfe01;
			16'hf281: y = 16'hfe01;
			16'hf282: y = 16'hfe01;
			16'hf283: y = 16'hfe01;
			16'hf284: y = 16'hfe01;
			16'hf285: y = 16'hfe01;
			16'hf286: y = 16'hfe01;
			16'hf287: y = 16'hfe01;
			16'hf288: y = 16'hfe01;
			16'hf289: y = 16'hfe01;
			16'hf28a: y = 16'hfe01;
			16'hf28b: y = 16'hfe01;
			16'hf28c: y = 16'hfe01;
			16'hf28d: y = 16'hfe01;
			16'hf28e: y = 16'hfe01;
			16'hf28f: y = 16'hfe01;
			16'hf290: y = 16'hfe01;
			16'hf291: y = 16'hfe01;
			16'hf292: y = 16'hfe01;
			16'hf293: y = 16'hfe01;
			16'hf294: y = 16'hfe01;
			16'hf295: y = 16'hfe01;
			16'hf296: y = 16'hfe01;
			16'hf297: y = 16'hfe01;
			16'hf298: y = 16'hfe01;
			16'hf299: y = 16'hfe01;
			16'hf29a: y = 16'hfe01;
			16'hf29b: y = 16'hfe01;
			16'hf29c: y = 16'hfe01;
			16'hf29d: y = 16'hfe01;
			16'hf29e: y = 16'hfe01;
			16'hf29f: y = 16'hfe01;
			16'hf2a0: y = 16'hfe01;
			16'hf2a1: y = 16'hfe01;
			16'hf2a2: y = 16'hfe01;
			16'hf2a3: y = 16'hfe01;
			16'hf2a4: y = 16'hfe01;
			16'hf2a5: y = 16'hfe01;
			16'hf2a6: y = 16'hfe01;
			16'hf2a7: y = 16'hfe01;
			16'hf2a8: y = 16'hfe01;
			16'hf2a9: y = 16'hfe01;
			16'hf2aa: y = 16'hfe01;
			16'hf2ab: y = 16'hfe01;
			16'hf2ac: y = 16'hfe01;
			16'hf2ad: y = 16'hfe01;
			16'hf2ae: y = 16'hfe01;
			16'hf2af: y = 16'hfe01;
			16'hf2b0: y = 16'hfe01;
			16'hf2b1: y = 16'hfe01;
			16'hf2b2: y = 16'hfe01;
			16'hf2b3: y = 16'hfe01;
			16'hf2b4: y = 16'hfe01;
			16'hf2b5: y = 16'hfe01;
			16'hf2b6: y = 16'hfe01;
			16'hf2b7: y = 16'hfe01;
			16'hf2b8: y = 16'hfe01;
			16'hf2b9: y = 16'hfe01;
			16'hf2ba: y = 16'hfe01;
			16'hf2bb: y = 16'hfe01;
			16'hf2bc: y = 16'hfe01;
			16'hf2bd: y = 16'hfe01;
			16'hf2be: y = 16'hfe01;
			16'hf2bf: y = 16'hfe01;
			16'hf2c0: y = 16'hfe01;
			16'hf2c1: y = 16'hfe01;
			16'hf2c2: y = 16'hfe01;
			16'hf2c3: y = 16'hfe01;
			16'hf2c4: y = 16'hfe01;
			16'hf2c5: y = 16'hfe01;
			16'hf2c6: y = 16'hfe01;
			16'hf2c7: y = 16'hfe01;
			16'hf2c8: y = 16'hfe01;
			16'hf2c9: y = 16'hfe01;
			16'hf2ca: y = 16'hfe01;
			16'hf2cb: y = 16'hfe01;
			16'hf2cc: y = 16'hfe01;
			16'hf2cd: y = 16'hfe01;
			16'hf2ce: y = 16'hfe01;
			16'hf2cf: y = 16'hfe01;
			16'hf2d0: y = 16'hfe01;
			16'hf2d1: y = 16'hfe01;
			16'hf2d2: y = 16'hfe01;
			16'hf2d3: y = 16'hfe01;
			16'hf2d4: y = 16'hfe01;
			16'hf2d5: y = 16'hfe01;
			16'hf2d6: y = 16'hfe01;
			16'hf2d7: y = 16'hfe01;
			16'hf2d8: y = 16'hfe01;
			16'hf2d9: y = 16'hfe01;
			16'hf2da: y = 16'hfe01;
			16'hf2db: y = 16'hfe01;
			16'hf2dc: y = 16'hfe01;
			16'hf2dd: y = 16'hfe01;
			16'hf2de: y = 16'hfe01;
			16'hf2df: y = 16'hfe01;
			16'hf2e0: y = 16'hfe01;
			16'hf2e1: y = 16'hfe01;
			16'hf2e2: y = 16'hfe01;
			16'hf2e3: y = 16'hfe01;
			16'hf2e4: y = 16'hfe01;
			16'hf2e5: y = 16'hfe01;
			16'hf2e6: y = 16'hfe01;
			16'hf2e7: y = 16'hfe01;
			16'hf2e8: y = 16'hfe01;
			16'hf2e9: y = 16'hfe01;
			16'hf2ea: y = 16'hfe01;
			16'hf2eb: y = 16'hfe01;
			16'hf2ec: y = 16'hfe01;
			16'hf2ed: y = 16'hfe01;
			16'hf2ee: y = 16'hfe01;
			16'hf2ef: y = 16'hfe01;
			16'hf2f0: y = 16'hfe01;
			16'hf2f1: y = 16'hfe01;
			16'hf2f2: y = 16'hfe01;
			16'hf2f3: y = 16'hfe01;
			16'hf2f4: y = 16'hfe01;
			16'hf2f5: y = 16'hfe01;
			16'hf2f6: y = 16'hfe01;
			16'hf2f7: y = 16'hfe01;
			16'hf2f8: y = 16'hfe01;
			16'hf2f9: y = 16'hfe01;
			16'hf2fa: y = 16'hfe01;
			16'hf2fb: y = 16'hfe01;
			16'hf2fc: y = 16'hfe01;
			16'hf2fd: y = 16'hfe01;
			16'hf2fe: y = 16'hfe01;
			16'hf2ff: y = 16'hfe01;
			16'hf300: y = 16'hfe01;
			16'hf301: y = 16'hfe01;
			16'hf302: y = 16'hfe01;
			16'hf303: y = 16'hfe01;
			16'hf304: y = 16'hfe01;
			16'hf305: y = 16'hfe01;
			16'hf306: y = 16'hfe01;
			16'hf307: y = 16'hfe01;
			16'hf308: y = 16'hfe01;
			16'hf309: y = 16'hfe01;
			16'hf30a: y = 16'hfe01;
			16'hf30b: y = 16'hfe01;
			16'hf30c: y = 16'hfe01;
			16'hf30d: y = 16'hfe01;
			16'hf30e: y = 16'hfe01;
			16'hf30f: y = 16'hfe01;
			16'hf310: y = 16'hfe01;
			16'hf311: y = 16'hfe01;
			16'hf312: y = 16'hfe01;
			16'hf313: y = 16'hfe01;
			16'hf314: y = 16'hfe01;
			16'hf315: y = 16'hfe01;
			16'hf316: y = 16'hfe01;
			16'hf317: y = 16'hfe01;
			16'hf318: y = 16'hfe01;
			16'hf319: y = 16'hfe01;
			16'hf31a: y = 16'hfe01;
			16'hf31b: y = 16'hfe01;
			16'hf31c: y = 16'hfe01;
			16'hf31d: y = 16'hfe01;
			16'hf31e: y = 16'hfe01;
			16'hf31f: y = 16'hfe01;
			16'hf320: y = 16'hfe01;
			16'hf321: y = 16'hfe01;
			16'hf322: y = 16'hfe01;
			16'hf323: y = 16'hfe01;
			16'hf324: y = 16'hfe01;
			16'hf325: y = 16'hfe01;
			16'hf326: y = 16'hfe01;
			16'hf327: y = 16'hfe01;
			16'hf328: y = 16'hfe01;
			16'hf329: y = 16'hfe01;
			16'hf32a: y = 16'hfe01;
			16'hf32b: y = 16'hfe01;
			16'hf32c: y = 16'hfe01;
			16'hf32d: y = 16'hfe01;
			16'hf32e: y = 16'hfe01;
			16'hf32f: y = 16'hfe01;
			16'hf330: y = 16'hfe01;
			16'hf331: y = 16'hfe01;
			16'hf332: y = 16'hfe01;
			16'hf333: y = 16'hfe01;
			16'hf334: y = 16'hfe01;
			16'hf335: y = 16'hfe01;
			16'hf336: y = 16'hfe01;
			16'hf337: y = 16'hfe01;
			16'hf338: y = 16'hfe01;
			16'hf339: y = 16'hfe01;
			16'hf33a: y = 16'hfe01;
			16'hf33b: y = 16'hfe01;
			16'hf33c: y = 16'hfe01;
			16'hf33d: y = 16'hfe01;
			16'hf33e: y = 16'hfe01;
			16'hf33f: y = 16'hfe01;
			16'hf340: y = 16'hfe01;
			16'hf341: y = 16'hfe01;
			16'hf342: y = 16'hfe01;
			16'hf343: y = 16'hfe01;
			16'hf344: y = 16'hfe01;
			16'hf345: y = 16'hfe01;
			16'hf346: y = 16'hfe01;
			16'hf347: y = 16'hfe01;
			16'hf348: y = 16'hfe01;
			16'hf349: y = 16'hfe01;
			16'hf34a: y = 16'hfe01;
			16'hf34b: y = 16'hfe01;
			16'hf34c: y = 16'hfe01;
			16'hf34d: y = 16'hfe01;
			16'hf34e: y = 16'hfe01;
			16'hf34f: y = 16'hfe01;
			16'hf350: y = 16'hfe01;
			16'hf351: y = 16'hfe01;
			16'hf352: y = 16'hfe01;
			16'hf353: y = 16'hfe01;
			16'hf354: y = 16'hfe01;
			16'hf355: y = 16'hfe01;
			16'hf356: y = 16'hfe01;
			16'hf357: y = 16'hfe01;
			16'hf358: y = 16'hfe01;
			16'hf359: y = 16'hfe01;
			16'hf35a: y = 16'hfe01;
			16'hf35b: y = 16'hfe01;
			16'hf35c: y = 16'hfe01;
			16'hf35d: y = 16'hfe01;
			16'hf35e: y = 16'hfe01;
			16'hf35f: y = 16'hfe01;
			16'hf360: y = 16'hfe01;
			16'hf361: y = 16'hfe01;
			16'hf362: y = 16'hfe01;
			16'hf363: y = 16'hfe01;
			16'hf364: y = 16'hfe01;
			16'hf365: y = 16'hfe01;
			16'hf366: y = 16'hfe01;
			16'hf367: y = 16'hfe01;
			16'hf368: y = 16'hfe01;
			16'hf369: y = 16'hfe01;
			16'hf36a: y = 16'hfe01;
			16'hf36b: y = 16'hfe01;
			16'hf36c: y = 16'hfe01;
			16'hf36d: y = 16'hfe01;
			16'hf36e: y = 16'hfe01;
			16'hf36f: y = 16'hfe01;
			16'hf370: y = 16'hfe01;
			16'hf371: y = 16'hfe01;
			16'hf372: y = 16'hfe01;
			16'hf373: y = 16'hfe01;
			16'hf374: y = 16'hfe01;
			16'hf375: y = 16'hfe01;
			16'hf376: y = 16'hfe01;
			16'hf377: y = 16'hfe01;
			16'hf378: y = 16'hfe01;
			16'hf379: y = 16'hfe01;
			16'hf37a: y = 16'hfe01;
			16'hf37b: y = 16'hfe01;
			16'hf37c: y = 16'hfe01;
			16'hf37d: y = 16'hfe01;
			16'hf37e: y = 16'hfe01;
			16'hf37f: y = 16'hfe01;
			16'hf380: y = 16'hfe01;
			16'hf381: y = 16'hfe01;
			16'hf382: y = 16'hfe01;
			16'hf383: y = 16'hfe01;
			16'hf384: y = 16'hfe01;
			16'hf385: y = 16'hfe01;
			16'hf386: y = 16'hfe01;
			16'hf387: y = 16'hfe01;
			16'hf388: y = 16'hfe01;
			16'hf389: y = 16'hfe01;
			16'hf38a: y = 16'hfe01;
			16'hf38b: y = 16'hfe01;
			16'hf38c: y = 16'hfe01;
			16'hf38d: y = 16'hfe01;
			16'hf38e: y = 16'hfe01;
			16'hf38f: y = 16'hfe01;
			16'hf390: y = 16'hfe01;
			16'hf391: y = 16'hfe01;
			16'hf392: y = 16'hfe01;
			16'hf393: y = 16'hfe01;
			16'hf394: y = 16'hfe01;
			16'hf395: y = 16'hfe01;
			16'hf396: y = 16'hfe01;
			16'hf397: y = 16'hfe01;
			16'hf398: y = 16'hfe01;
			16'hf399: y = 16'hfe01;
			16'hf39a: y = 16'hfe01;
			16'hf39b: y = 16'hfe01;
			16'hf39c: y = 16'hfe01;
			16'hf39d: y = 16'hfe01;
			16'hf39e: y = 16'hfe01;
			16'hf39f: y = 16'hfe01;
			16'hf3a0: y = 16'hfe01;
			16'hf3a1: y = 16'hfe01;
			16'hf3a2: y = 16'hfe01;
			16'hf3a3: y = 16'hfe01;
			16'hf3a4: y = 16'hfe01;
			16'hf3a5: y = 16'hfe01;
			16'hf3a6: y = 16'hfe01;
			16'hf3a7: y = 16'hfe01;
			16'hf3a8: y = 16'hfe01;
			16'hf3a9: y = 16'hfe01;
			16'hf3aa: y = 16'hfe01;
			16'hf3ab: y = 16'hfe01;
			16'hf3ac: y = 16'hfe01;
			16'hf3ad: y = 16'hfe01;
			16'hf3ae: y = 16'hfe01;
			16'hf3af: y = 16'hfe01;
			16'hf3b0: y = 16'hfe01;
			16'hf3b1: y = 16'hfe01;
			16'hf3b2: y = 16'hfe01;
			16'hf3b3: y = 16'hfe01;
			16'hf3b4: y = 16'hfe01;
			16'hf3b5: y = 16'hfe01;
			16'hf3b6: y = 16'hfe01;
			16'hf3b7: y = 16'hfe01;
			16'hf3b8: y = 16'hfe01;
			16'hf3b9: y = 16'hfe01;
			16'hf3ba: y = 16'hfe01;
			16'hf3bb: y = 16'hfe01;
			16'hf3bc: y = 16'hfe01;
			16'hf3bd: y = 16'hfe01;
			16'hf3be: y = 16'hfe01;
			16'hf3bf: y = 16'hfe01;
			16'hf3c0: y = 16'hfe01;
			16'hf3c1: y = 16'hfe01;
			16'hf3c2: y = 16'hfe01;
			16'hf3c3: y = 16'hfe01;
			16'hf3c4: y = 16'hfe01;
			16'hf3c5: y = 16'hfe01;
			16'hf3c6: y = 16'hfe01;
			16'hf3c7: y = 16'hfe01;
			16'hf3c8: y = 16'hfe01;
			16'hf3c9: y = 16'hfe01;
			16'hf3ca: y = 16'hfe01;
			16'hf3cb: y = 16'hfe01;
			16'hf3cc: y = 16'hfe01;
			16'hf3cd: y = 16'hfe01;
			16'hf3ce: y = 16'hfe01;
			16'hf3cf: y = 16'hfe01;
			16'hf3d0: y = 16'hfe01;
			16'hf3d1: y = 16'hfe01;
			16'hf3d2: y = 16'hfe01;
			16'hf3d3: y = 16'hfe01;
			16'hf3d4: y = 16'hfe01;
			16'hf3d5: y = 16'hfe01;
			16'hf3d6: y = 16'hfe01;
			16'hf3d7: y = 16'hfe01;
			16'hf3d8: y = 16'hfe01;
			16'hf3d9: y = 16'hfe01;
			16'hf3da: y = 16'hfe01;
			16'hf3db: y = 16'hfe01;
			16'hf3dc: y = 16'hfe01;
			16'hf3dd: y = 16'hfe01;
			16'hf3de: y = 16'hfe01;
			16'hf3df: y = 16'hfe01;
			16'hf3e0: y = 16'hfe01;
			16'hf3e1: y = 16'hfe01;
			16'hf3e2: y = 16'hfe01;
			16'hf3e3: y = 16'hfe01;
			16'hf3e4: y = 16'hfe01;
			16'hf3e5: y = 16'hfe01;
			16'hf3e6: y = 16'hfe01;
			16'hf3e7: y = 16'hfe01;
			16'hf3e8: y = 16'hfe01;
			16'hf3e9: y = 16'hfe01;
			16'hf3ea: y = 16'hfe01;
			16'hf3eb: y = 16'hfe01;
			16'hf3ec: y = 16'hfe01;
			16'hf3ed: y = 16'hfe01;
			16'hf3ee: y = 16'hfe01;
			16'hf3ef: y = 16'hfe01;
			16'hf3f0: y = 16'hfe01;
			16'hf3f1: y = 16'hfe01;
			16'hf3f2: y = 16'hfe01;
			16'hf3f3: y = 16'hfe01;
			16'hf3f4: y = 16'hfe01;
			16'hf3f5: y = 16'hfe01;
			16'hf3f6: y = 16'hfe01;
			16'hf3f7: y = 16'hfe01;
			16'hf3f8: y = 16'hfe01;
			16'hf3f9: y = 16'hfe01;
			16'hf3fa: y = 16'hfe01;
			16'hf3fb: y = 16'hfe01;
			16'hf3fc: y = 16'hfe01;
			16'hf3fd: y = 16'hfe01;
			16'hf3fe: y = 16'hfe01;
			16'hf3ff: y = 16'hfe01;
			16'hf400: y = 16'hfe01;
			16'hf401: y = 16'hfe01;
			16'hf402: y = 16'hfe01;
			16'hf403: y = 16'hfe01;
			16'hf404: y = 16'hfe01;
			16'hf405: y = 16'hfe01;
			16'hf406: y = 16'hfe01;
			16'hf407: y = 16'hfe01;
			16'hf408: y = 16'hfe01;
			16'hf409: y = 16'hfe01;
			16'hf40a: y = 16'hfe01;
			16'hf40b: y = 16'hfe01;
			16'hf40c: y = 16'hfe01;
			16'hf40d: y = 16'hfe01;
			16'hf40e: y = 16'hfe01;
			16'hf40f: y = 16'hfe01;
			16'hf410: y = 16'hfe01;
			16'hf411: y = 16'hfe01;
			16'hf412: y = 16'hfe01;
			16'hf413: y = 16'hfe01;
			16'hf414: y = 16'hfe01;
			16'hf415: y = 16'hfe01;
			16'hf416: y = 16'hfe01;
			16'hf417: y = 16'hfe01;
			16'hf418: y = 16'hfe01;
			16'hf419: y = 16'hfe01;
			16'hf41a: y = 16'hfe01;
			16'hf41b: y = 16'hfe01;
			16'hf41c: y = 16'hfe01;
			16'hf41d: y = 16'hfe01;
			16'hf41e: y = 16'hfe01;
			16'hf41f: y = 16'hfe01;
			16'hf420: y = 16'hfe01;
			16'hf421: y = 16'hfe01;
			16'hf422: y = 16'hfe01;
			16'hf423: y = 16'hfe01;
			16'hf424: y = 16'hfe01;
			16'hf425: y = 16'hfe01;
			16'hf426: y = 16'hfe01;
			16'hf427: y = 16'hfe01;
			16'hf428: y = 16'hfe01;
			16'hf429: y = 16'hfe01;
			16'hf42a: y = 16'hfe01;
			16'hf42b: y = 16'hfe01;
			16'hf42c: y = 16'hfe01;
			16'hf42d: y = 16'hfe01;
			16'hf42e: y = 16'hfe01;
			16'hf42f: y = 16'hfe01;
			16'hf430: y = 16'hfe01;
			16'hf431: y = 16'hfe01;
			16'hf432: y = 16'hfe01;
			16'hf433: y = 16'hfe01;
			16'hf434: y = 16'hfe01;
			16'hf435: y = 16'hfe01;
			16'hf436: y = 16'hfe01;
			16'hf437: y = 16'hfe01;
			16'hf438: y = 16'hfe01;
			16'hf439: y = 16'hfe01;
			16'hf43a: y = 16'hfe01;
			16'hf43b: y = 16'hfe01;
			16'hf43c: y = 16'hfe01;
			16'hf43d: y = 16'hfe01;
			16'hf43e: y = 16'hfe01;
			16'hf43f: y = 16'hfe01;
			16'hf440: y = 16'hfe01;
			16'hf441: y = 16'hfe01;
			16'hf442: y = 16'hfe01;
			16'hf443: y = 16'hfe01;
			16'hf444: y = 16'hfe01;
			16'hf445: y = 16'hfe01;
			16'hf446: y = 16'hfe01;
			16'hf447: y = 16'hfe01;
			16'hf448: y = 16'hfe01;
			16'hf449: y = 16'hfe01;
			16'hf44a: y = 16'hfe01;
			16'hf44b: y = 16'hfe01;
			16'hf44c: y = 16'hfe01;
			16'hf44d: y = 16'hfe01;
			16'hf44e: y = 16'hfe01;
			16'hf44f: y = 16'hfe01;
			16'hf450: y = 16'hfe01;
			16'hf451: y = 16'hfe01;
			16'hf452: y = 16'hfe01;
			16'hf453: y = 16'hfe01;
			16'hf454: y = 16'hfe01;
			16'hf455: y = 16'hfe01;
			16'hf456: y = 16'hfe01;
			16'hf457: y = 16'hfe01;
			16'hf458: y = 16'hfe01;
			16'hf459: y = 16'hfe01;
			16'hf45a: y = 16'hfe01;
			16'hf45b: y = 16'hfe01;
			16'hf45c: y = 16'hfe01;
			16'hf45d: y = 16'hfe01;
			16'hf45e: y = 16'hfe01;
			16'hf45f: y = 16'hfe01;
			16'hf460: y = 16'hfe01;
			16'hf461: y = 16'hfe01;
			16'hf462: y = 16'hfe01;
			16'hf463: y = 16'hfe01;
			16'hf464: y = 16'hfe01;
			16'hf465: y = 16'hfe01;
			16'hf466: y = 16'hfe01;
			16'hf467: y = 16'hfe01;
			16'hf468: y = 16'hfe01;
			16'hf469: y = 16'hfe01;
			16'hf46a: y = 16'hfe01;
			16'hf46b: y = 16'hfe01;
			16'hf46c: y = 16'hfe01;
			16'hf46d: y = 16'hfe01;
			16'hf46e: y = 16'hfe01;
			16'hf46f: y = 16'hfe01;
			16'hf470: y = 16'hfe01;
			16'hf471: y = 16'hfe01;
			16'hf472: y = 16'hfe01;
			16'hf473: y = 16'hfe01;
			16'hf474: y = 16'hfe01;
			16'hf475: y = 16'hfe01;
			16'hf476: y = 16'hfe01;
			16'hf477: y = 16'hfe01;
			16'hf478: y = 16'hfe01;
			16'hf479: y = 16'hfe01;
			16'hf47a: y = 16'hfe01;
			16'hf47b: y = 16'hfe01;
			16'hf47c: y = 16'hfe01;
			16'hf47d: y = 16'hfe01;
			16'hf47e: y = 16'hfe01;
			16'hf47f: y = 16'hfe01;
			16'hf480: y = 16'hfe01;
			16'hf481: y = 16'hfe01;
			16'hf482: y = 16'hfe01;
			16'hf483: y = 16'hfe01;
			16'hf484: y = 16'hfe01;
			16'hf485: y = 16'hfe01;
			16'hf486: y = 16'hfe01;
			16'hf487: y = 16'hfe01;
			16'hf488: y = 16'hfe01;
			16'hf489: y = 16'hfe01;
			16'hf48a: y = 16'hfe01;
			16'hf48b: y = 16'hfe01;
			16'hf48c: y = 16'hfe01;
			16'hf48d: y = 16'hfe01;
			16'hf48e: y = 16'hfe01;
			16'hf48f: y = 16'hfe01;
			16'hf490: y = 16'hfe01;
			16'hf491: y = 16'hfe01;
			16'hf492: y = 16'hfe01;
			16'hf493: y = 16'hfe01;
			16'hf494: y = 16'hfe01;
			16'hf495: y = 16'hfe01;
			16'hf496: y = 16'hfe01;
			16'hf497: y = 16'hfe01;
			16'hf498: y = 16'hfe01;
			16'hf499: y = 16'hfe01;
			16'hf49a: y = 16'hfe01;
			16'hf49b: y = 16'hfe01;
			16'hf49c: y = 16'hfe01;
			16'hf49d: y = 16'hfe01;
			16'hf49e: y = 16'hfe01;
			16'hf49f: y = 16'hfe01;
			16'hf4a0: y = 16'hfe01;
			16'hf4a1: y = 16'hfe01;
			16'hf4a2: y = 16'hfe01;
			16'hf4a3: y = 16'hfe01;
			16'hf4a4: y = 16'hfe01;
			16'hf4a5: y = 16'hfe01;
			16'hf4a6: y = 16'hfe01;
			16'hf4a7: y = 16'hfe01;
			16'hf4a8: y = 16'hfe01;
			16'hf4a9: y = 16'hfe01;
			16'hf4aa: y = 16'hfe01;
			16'hf4ab: y = 16'hfe01;
			16'hf4ac: y = 16'hfe01;
			16'hf4ad: y = 16'hfe01;
			16'hf4ae: y = 16'hfe01;
			16'hf4af: y = 16'hfe01;
			16'hf4b0: y = 16'hfe01;
			16'hf4b1: y = 16'hfe01;
			16'hf4b2: y = 16'hfe01;
			16'hf4b3: y = 16'hfe01;
			16'hf4b4: y = 16'hfe01;
			16'hf4b5: y = 16'hfe01;
			16'hf4b6: y = 16'hfe01;
			16'hf4b7: y = 16'hfe01;
			16'hf4b8: y = 16'hfe01;
			16'hf4b9: y = 16'hfe01;
			16'hf4ba: y = 16'hfe01;
			16'hf4bb: y = 16'hfe01;
			16'hf4bc: y = 16'hfe01;
			16'hf4bd: y = 16'hfe01;
			16'hf4be: y = 16'hfe01;
			16'hf4bf: y = 16'hfe01;
			16'hf4c0: y = 16'hfe01;
			16'hf4c1: y = 16'hfe01;
			16'hf4c2: y = 16'hfe01;
			16'hf4c3: y = 16'hfe01;
			16'hf4c4: y = 16'hfe01;
			16'hf4c5: y = 16'hfe01;
			16'hf4c6: y = 16'hfe01;
			16'hf4c7: y = 16'hfe01;
			16'hf4c8: y = 16'hfe01;
			16'hf4c9: y = 16'hfe01;
			16'hf4ca: y = 16'hfe01;
			16'hf4cb: y = 16'hfe01;
			16'hf4cc: y = 16'hfe01;
			16'hf4cd: y = 16'hfe01;
			16'hf4ce: y = 16'hfe01;
			16'hf4cf: y = 16'hfe01;
			16'hf4d0: y = 16'hfe01;
			16'hf4d1: y = 16'hfe01;
			16'hf4d2: y = 16'hfe01;
			16'hf4d3: y = 16'hfe01;
			16'hf4d4: y = 16'hfe01;
			16'hf4d5: y = 16'hfe01;
			16'hf4d6: y = 16'hfe01;
			16'hf4d7: y = 16'hfe01;
			16'hf4d8: y = 16'hfe01;
			16'hf4d9: y = 16'hfe01;
			16'hf4da: y = 16'hfe01;
			16'hf4db: y = 16'hfe01;
			16'hf4dc: y = 16'hfe01;
			16'hf4dd: y = 16'hfe01;
			16'hf4de: y = 16'hfe01;
			16'hf4df: y = 16'hfe01;
			16'hf4e0: y = 16'hfe01;
			16'hf4e1: y = 16'hfe01;
			16'hf4e2: y = 16'hfe01;
			16'hf4e3: y = 16'hfe01;
			16'hf4e4: y = 16'hfe01;
			16'hf4e5: y = 16'hfe01;
			16'hf4e6: y = 16'hfe01;
			16'hf4e7: y = 16'hfe01;
			16'hf4e8: y = 16'hfe01;
			16'hf4e9: y = 16'hfe01;
			16'hf4ea: y = 16'hfe01;
			16'hf4eb: y = 16'hfe01;
			16'hf4ec: y = 16'hfe01;
			16'hf4ed: y = 16'hfe01;
			16'hf4ee: y = 16'hfe01;
			16'hf4ef: y = 16'hfe01;
			16'hf4f0: y = 16'hfe01;
			16'hf4f1: y = 16'hfe01;
			16'hf4f2: y = 16'hfe01;
			16'hf4f3: y = 16'hfe01;
			16'hf4f4: y = 16'hfe01;
			16'hf4f5: y = 16'hfe01;
			16'hf4f6: y = 16'hfe01;
			16'hf4f7: y = 16'hfe01;
			16'hf4f8: y = 16'hfe01;
			16'hf4f9: y = 16'hfe01;
			16'hf4fa: y = 16'hfe01;
			16'hf4fb: y = 16'hfe01;
			16'hf4fc: y = 16'hfe01;
			16'hf4fd: y = 16'hfe01;
			16'hf4fe: y = 16'hfe01;
			16'hf4ff: y = 16'hfe01;
			16'hf500: y = 16'hfe01;
			16'hf501: y = 16'hfe01;
			16'hf502: y = 16'hfe01;
			16'hf503: y = 16'hfe01;
			16'hf504: y = 16'hfe01;
			16'hf505: y = 16'hfe01;
			16'hf506: y = 16'hfe01;
			16'hf507: y = 16'hfe01;
			16'hf508: y = 16'hfe01;
			16'hf509: y = 16'hfe01;
			16'hf50a: y = 16'hfe01;
			16'hf50b: y = 16'hfe01;
			16'hf50c: y = 16'hfe01;
			16'hf50d: y = 16'hfe01;
			16'hf50e: y = 16'hfe01;
			16'hf50f: y = 16'hfe01;
			16'hf510: y = 16'hfe01;
			16'hf511: y = 16'hfe01;
			16'hf512: y = 16'hfe01;
			16'hf513: y = 16'hfe01;
			16'hf514: y = 16'hfe01;
			16'hf515: y = 16'hfe01;
			16'hf516: y = 16'hfe01;
			16'hf517: y = 16'hfe01;
			16'hf518: y = 16'hfe01;
			16'hf519: y = 16'hfe01;
			16'hf51a: y = 16'hfe01;
			16'hf51b: y = 16'hfe01;
			16'hf51c: y = 16'hfe01;
			16'hf51d: y = 16'hfe01;
			16'hf51e: y = 16'hfe01;
			16'hf51f: y = 16'hfe01;
			16'hf520: y = 16'hfe01;
			16'hf521: y = 16'hfe01;
			16'hf522: y = 16'hfe01;
			16'hf523: y = 16'hfe01;
			16'hf524: y = 16'hfe01;
			16'hf525: y = 16'hfe01;
			16'hf526: y = 16'hfe01;
			16'hf527: y = 16'hfe01;
			16'hf528: y = 16'hfe01;
			16'hf529: y = 16'hfe01;
			16'hf52a: y = 16'hfe01;
			16'hf52b: y = 16'hfe01;
			16'hf52c: y = 16'hfe01;
			16'hf52d: y = 16'hfe01;
			16'hf52e: y = 16'hfe01;
			16'hf52f: y = 16'hfe01;
			16'hf530: y = 16'hfe01;
			16'hf531: y = 16'hfe01;
			16'hf532: y = 16'hfe01;
			16'hf533: y = 16'hfe01;
			16'hf534: y = 16'hfe01;
			16'hf535: y = 16'hfe01;
			16'hf536: y = 16'hfe01;
			16'hf537: y = 16'hfe01;
			16'hf538: y = 16'hfe01;
			16'hf539: y = 16'hfe01;
			16'hf53a: y = 16'hfe01;
			16'hf53b: y = 16'hfe01;
			16'hf53c: y = 16'hfe01;
			16'hf53d: y = 16'hfe01;
			16'hf53e: y = 16'hfe01;
			16'hf53f: y = 16'hfe01;
			16'hf540: y = 16'hfe01;
			16'hf541: y = 16'hfe01;
			16'hf542: y = 16'hfe01;
			16'hf543: y = 16'hfe01;
			16'hf544: y = 16'hfe01;
			16'hf545: y = 16'hfe01;
			16'hf546: y = 16'hfe01;
			16'hf547: y = 16'hfe01;
			16'hf548: y = 16'hfe01;
			16'hf549: y = 16'hfe01;
			16'hf54a: y = 16'hfe01;
			16'hf54b: y = 16'hfe01;
			16'hf54c: y = 16'hfe01;
			16'hf54d: y = 16'hfe01;
			16'hf54e: y = 16'hfe01;
			16'hf54f: y = 16'hfe01;
			16'hf550: y = 16'hfe01;
			16'hf551: y = 16'hfe01;
			16'hf552: y = 16'hfe01;
			16'hf553: y = 16'hfe01;
			16'hf554: y = 16'hfe01;
			16'hf555: y = 16'hfe01;
			16'hf556: y = 16'hfe01;
			16'hf557: y = 16'hfe01;
			16'hf558: y = 16'hfe01;
			16'hf559: y = 16'hfe01;
			16'hf55a: y = 16'hfe01;
			16'hf55b: y = 16'hfe01;
			16'hf55c: y = 16'hfe01;
			16'hf55d: y = 16'hfe01;
			16'hf55e: y = 16'hfe01;
			16'hf55f: y = 16'hfe01;
			16'hf560: y = 16'hfe01;
			16'hf561: y = 16'hfe01;
			16'hf562: y = 16'hfe01;
			16'hf563: y = 16'hfe01;
			16'hf564: y = 16'hfe01;
			16'hf565: y = 16'hfe01;
			16'hf566: y = 16'hfe01;
			16'hf567: y = 16'hfe01;
			16'hf568: y = 16'hfe01;
			16'hf569: y = 16'hfe01;
			16'hf56a: y = 16'hfe01;
			16'hf56b: y = 16'hfe01;
			16'hf56c: y = 16'hfe01;
			16'hf56d: y = 16'hfe01;
			16'hf56e: y = 16'hfe01;
			16'hf56f: y = 16'hfe01;
			16'hf570: y = 16'hfe01;
			16'hf571: y = 16'hfe01;
			16'hf572: y = 16'hfe01;
			16'hf573: y = 16'hfe01;
			16'hf574: y = 16'hfe01;
			16'hf575: y = 16'hfe01;
			16'hf576: y = 16'hfe01;
			16'hf577: y = 16'hfe01;
			16'hf578: y = 16'hfe01;
			16'hf579: y = 16'hfe01;
			16'hf57a: y = 16'hfe01;
			16'hf57b: y = 16'hfe01;
			16'hf57c: y = 16'hfe01;
			16'hf57d: y = 16'hfe01;
			16'hf57e: y = 16'hfe01;
			16'hf57f: y = 16'hfe01;
			16'hf580: y = 16'hfe01;
			16'hf581: y = 16'hfe01;
			16'hf582: y = 16'hfe01;
			16'hf583: y = 16'hfe01;
			16'hf584: y = 16'hfe01;
			16'hf585: y = 16'hfe01;
			16'hf586: y = 16'hfe01;
			16'hf587: y = 16'hfe01;
			16'hf588: y = 16'hfe01;
			16'hf589: y = 16'hfe01;
			16'hf58a: y = 16'hfe01;
			16'hf58b: y = 16'hfe01;
			16'hf58c: y = 16'hfe01;
			16'hf58d: y = 16'hfe01;
			16'hf58e: y = 16'hfe01;
			16'hf58f: y = 16'hfe01;
			16'hf590: y = 16'hfe01;
			16'hf591: y = 16'hfe01;
			16'hf592: y = 16'hfe01;
			16'hf593: y = 16'hfe01;
			16'hf594: y = 16'hfe01;
			16'hf595: y = 16'hfe01;
			16'hf596: y = 16'hfe01;
			16'hf597: y = 16'hfe01;
			16'hf598: y = 16'hfe01;
			16'hf599: y = 16'hfe01;
			16'hf59a: y = 16'hfe01;
			16'hf59b: y = 16'hfe01;
			16'hf59c: y = 16'hfe01;
			16'hf59d: y = 16'hfe01;
			16'hf59e: y = 16'hfe01;
			16'hf59f: y = 16'hfe01;
			16'hf5a0: y = 16'hfe01;
			16'hf5a1: y = 16'hfe01;
			16'hf5a2: y = 16'hfe01;
			16'hf5a3: y = 16'hfe01;
			16'hf5a4: y = 16'hfe01;
			16'hf5a5: y = 16'hfe01;
			16'hf5a6: y = 16'hfe01;
			16'hf5a7: y = 16'hfe01;
			16'hf5a8: y = 16'hfe01;
			16'hf5a9: y = 16'hfe01;
			16'hf5aa: y = 16'hfe01;
			16'hf5ab: y = 16'hfe01;
			16'hf5ac: y = 16'hfe01;
			16'hf5ad: y = 16'hfe01;
			16'hf5ae: y = 16'hfe01;
			16'hf5af: y = 16'hfe01;
			16'hf5b0: y = 16'hfe01;
			16'hf5b1: y = 16'hfe01;
			16'hf5b2: y = 16'hfe01;
			16'hf5b3: y = 16'hfe01;
			16'hf5b4: y = 16'hfe01;
			16'hf5b5: y = 16'hfe01;
			16'hf5b6: y = 16'hfe01;
			16'hf5b7: y = 16'hfe01;
			16'hf5b8: y = 16'hfe01;
			16'hf5b9: y = 16'hfe01;
			16'hf5ba: y = 16'hfe01;
			16'hf5bb: y = 16'hfe01;
			16'hf5bc: y = 16'hfe01;
			16'hf5bd: y = 16'hfe01;
			16'hf5be: y = 16'hfe01;
			16'hf5bf: y = 16'hfe01;
			16'hf5c0: y = 16'hfe01;
			16'hf5c1: y = 16'hfe01;
			16'hf5c2: y = 16'hfe01;
			16'hf5c3: y = 16'hfe01;
			16'hf5c4: y = 16'hfe01;
			16'hf5c5: y = 16'hfe01;
			16'hf5c6: y = 16'hfe01;
			16'hf5c7: y = 16'hfe01;
			16'hf5c8: y = 16'hfe01;
			16'hf5c9: y = 16'hfe01;
			16'hf5ca: y = 16'hfe01;
			16'hf5cb: y = 16'hfe01;
			16'hf5cc: y = 16'hfe01;
			16'hf5cd: y = 16'hfe01;
			16'hf5ce: y = 16'hfe01;
			16'hf5cf: y = 16'hfe01;
			16'hf5d0: y = 16'hfe01;
			16'hf5d1: y = 16'hfe01;
			16'hf5d2: y = 16'hfe01;
			16'hf5d3: y = 16'hfe01;
			16'hf5d4: y = 16'hfe01;
			16'hf5d5: y = 16'hfe01;
			16'hf5d6: y = 16'hfe01;
			16'hf5d7: y = 16'hfe01;
			16'hf5d8: y = 16'hfe01;
			16'hf5d9: y = 16'hfe01;
			16'hf5da: y = 16'hfe01;
			16'hf5db: y = 16'hfe01;
			16'hf5dc: y = 16'hfe01;
			16'hf5dd: y = 16'hfe01;
			16'hf5de: y = 16'hfe01;
			16'hf5df: y = 16'hfe01;
			16'hf5e0: y = 16'hfe01;
			16'hf5e1: y = 16'hfe01;
			16'hf5e2: y = 16'hfe01;
			16'hf5e3: y = 16'hfe01;
			16'hf5e4: y = 16'hfe01;
			16'hf5e5: y = 16'hfe01;
			16'hf5e6: y = 16'hfe01;
			16'hf5e7: y = 16'hfe01;
			16'hf5e8: y = 16'hfe01;
			16'hf5e9: y = 16'hfe01;
			16'hf5ea: y = 16'hfe01;
			16'hf5eb: y = 16'hfe01;
			16'hf5ec: y = 16'hfe01;
			16'hf5ed: y = 16'hfe01;
			16'hf5ee: y = 16'hfe01;
			16'hf5ef: y = 16'hfe01;
			16'hf5f0: y = 16'hfe01;
			16'hf5f1: y = 16'hfe01;
			16'hf5f2: y = 16'hfe01;
			16'hf5f3: y = 16'hfe01;
			16'hf5f4: y = 16'hfe01;
			16'hf5f5: y = 16'hfe01;
			16'hf5f6: y = 16'hfe01;
			16'hf5f7: y = 16'hfe01;
			16'hf5f8: y = 16'hfe01;
			16'hf5f9: y = 16'hfe01;
			16'hf5fa: y = 16'hfe01;
			16'hf5fb: y = 16'hfe01;
			16'hf5fc: y = 16'hfe01;
			16'hf5fd: y = 16'hfe01;
			16'hf5fe: y = 16'hfe01;
			16'hf5ff: y = 16'hfe01;
			16'hf600: y = 16'hfe01;
			16'hf601: y = 16'hfe01;
			16'hf602: y = 16'hfe01;
			16'hf603: y = 16'hfe01;
			16'hf604: y = 16'hfe01;
			16'hf605: y = 16'hfe01;
			16'hf606: y = 16'hfe01;
			16'hf607: y = 16'hfe01;
			16'hf608: y = 16'hfe01;
			16'hf609: y = 16'hfe01;
			16'hf60a: y = 16'hfe01;
			16'hf60b: y = 16'hfe01;
			16'hf60c: y = 16'hfe01;
			16'hf60d: y = 16'hfe01;
			16'hf60e: y = 16'hfe01;
			16'hf60f: y = 16'hfe01;
			16'hf610: y = 16'hfe01;
			16'hf611: y = 16'hfe01;
			16'hf612: y = 16'hfe01;
			16'hf613: y = 16'hfe01;
			16'hf614: y = 16'hfe01;
			16'hf615: y = 16'hfe01;
			16'hf616: y = 16'hfe01;
			16'hf617: y = 16'hfe01;
			16'hf618: y = 16'hfe01;
			16'hf619: y = 16'hfe01;
			16'hf61a: y = 16'hfe01;
			16'hf61b: y = 16'hfe01;
			16'hf61c: y = 16'hfe01;
			16'hf61d: y = 16'hfe01;
			16'hf61e: y = 16'hfe01;
			16'hf61f: y = 16'hfe01;
			16'hf620: y = 16'hfe01;
			16'hf621: y = 16'hfe01;
			16'hf622: y = 16'hfe01;
			16'hf623: y = 16'hfe01;
			16'hf624: y = 16'hfe01;
			16'hf625: y = 16'hfe01;
			16'hf626: y = 16'hfe01;
			16'hf627: y = 16'hfe01;
			16'hf628: y = 16'hfe01;
			16'hf629: y = 16'hfe01;
			16'hf62a: y = 16'hfe01;
			16'hf62b: y = 16'hfe01;
			16'hf62c: y = 16'hfe01;
			16'hf62d: y = 16'hfe01;
			16'hf62e: y = 16'hfe01;
			16'hf62f: y = 16'hfe01;
			16'hf630: y = 16'hfe01;
			16'hf631: y = 16'hfe01;
			16'hf632: y = 16'hfe01;
			16'hf633: y = 16'hfe01;
			16'hf634: y = 16'hfe01;
			16'hf635: y = 16'hfe01;
			16'hf636: y = 16'hfe01;
			16'hf637: y = 16'hfe01;
			16'hf638: y = 16'hfe01;
			16'hf639: y = 16'hfe01;
			16'hf63a: y = 16'hfe01;
			16'hf63b: y = 16'hfe01;
			16'hf63c: y = 16'hfe01;
			16'hf63d: y = 16'hfe01;
			16'hf63e: y = 16'hfe01;
			16'hf63f: y = 16'hfe01;
			16'hf640: y = 16'hfe01;
			16'hf641: y = 16'hfe01;
			16'hf642: y = 16'hfe01;
			16'hf643: y = 16'hfe01;
			16'hf644: y = 16'hfe01;
			16'hf645: y = 16'hfe01;
			16'hf646: y = 16'hfe01;
			16'hf647: y = 16'hfe01;
			16'hf648: y = 16'hfe01;
			16'hf649: y = 16'hfe01;
			16'hf64a: y = 16'hfe01;
			16'hf64b: y = 16'hfe01;
			16'hf64c: y = 16'hfe01;
			16'hf64d: y = 16'hfe01;
			16'hf64e: y = 16'hfe01;
			16'hf64f: y = 16'hfe01;
			16'hf650: y = 16'hfe01;
			16'hf651: y = 16'hfe01;
			16'hf652: y = 16'hfe01;
			16'hf653: y = 16'hfe01;
			16'hf654: y = 16'hfe01;
			16'hf655: y = 16'hfe01;
			16'hf656: y = 16'hfe01;
			16'hf657: y = 16'hfe01;
			16'hf658: y = 16'hfe01;
			16'hf659: y = 16'hfe01;
			16'hf65a: y = 16'hfe01;
			16'hf65b: y = 16'hfe01;
			16'hf65c: y = 16'hfe01;
			16'hf65d: y = 16'hfe01;
			16'hf65e: y = 16'hfe01;
			16'hf65f: y = 16'hfe01;
			16'hf660: y = 16'hfe01;
			16'hf661: y = 16'hfe01;
			16'hf662: y = 16'hfe01;
			16'hf663: y = 16'hfe01;
			16'hf664: y = 16'hfe01;
			16'hf665: y = 16'hfe01;
			16'hf666: y = 16'hfe01;
			16'hf667: y = 16'hfe01;
			16'hf668: y = 16'hfe01;
			16'hf669: y = 16'hfe01;
			16'hf66a: y = 16'hfe01;
			16'hf66b: y = 16'hfe01;
			16'hf66c: y = 16'hfe01;
			16'hf66d: y = 16'hfe01;
			16'hf66e: y = 16'hfe01;
			16'hf66f: y = 16'hfe01;
			16'hf670: y = 16'hfe01;
			16'hf671: y = 16'hfe01;
			16'hf672: y = 16'hfe01;
			16'hf673: y = 16'hfe01;
			16'hf674: y = 16'hfe01;
			16'hf675: y = 16'hfe01;
			16'hf676: y = 16'hfe01;
			16'hf677: y = 16'hfe01;
			16'hf678: y = 16'hfe01;
			16'hf679: y = 16'hfe01;
			16'hf67a: y = 16'hfe01;
			16'hf67b: y = 16'hfe01;
			16'hf67c: y = 16'hfe01;
			16'hf67d: y = 16'hfe01;
			16'hf67e: y = 16'hfe01;
			16'hf67f: y = 16'hfe01;
			16'hf680: y = 16'hfe01;
			16'hf681: y = 16'hfe01;
			16'hf682: y = 16'hfe01;
			16'hf683: y = 16'hfe01;
			16'hf684: y = 16'hfe01;
			16'hf685: y = 16'hfe01;
			16'hf686: y = 16'hfe01;
			16'hf687: y = 16'hfe01;
			16'hf688: y = 16'hfe01;
			16'hf689: y = 16'hfe01;
			16'hf68a: y = 16'hfe01;
			16'hf68b: y = 16'hfe01;
			16'hf68c: y = 16'hfe01;
			16'hf68d: y = 16'hfe01;
			16'hf68e: y = 16'hfe01;
			16'hf68f: y = 16'hfe01;
			16'hf690: y = 16'hfe01;
			16'hf691: y = 16'hfe01;
			16'hf692: y = 16'hfe01;
			16'hf693: y = 16'hfe01;
			16'hf694: y = 16'hfe01;
			16'hf695: y = 16'hfe01;
			16'hf696: y = 16'hfe01;
			16'hf697: y = 16'hfe01;
			16'hf698: y = 16'hfe01;
			16'hf699: y = 16'hfe01;
			16'hf69a: y = 16'hfe01;
			16'hf69b: y = 16'hfe01;
			16'hf69c: y = 16'hfe01;
			16'hf69d: y = 16'hfe01;
			16'hf69e: y = 16'hfe01;
			16'hf69f: y = 16'hfe01;
			16'hf6a0: y = 16'hfe01;
			16'hf6a1: y = 16'hfe01;
			16'hf6a2: y = 16'hfe01;
			16'hf6a3: y = 16'hfe01;
			16'hf6a4: y = 16'hfe01;
			16'hf6a5: y = 16'hfe01;
			16'hf6a6: y = 16'hfe01;
			16'hf6a7: y = 16'hfe01;
			16'hf6a8: y = 16'hfe01;
			16'hf6a9: y = 16'hfe01;
			16'hf6aa: y = 16'hfe01;
			16'hf6ab: y = 16'hfe01;
			16'hf6ac: y = 16'hfe01;
			16'hf6ad: y = 16'hfe01;
			16'hf6ae: y = 16'hfe01;
			16'hf6af: y = 16'hfe01;
			16'hf6b0: y = 16'hfe01;
			16'hf6b1: y = 16'hfe01;
			16'hf6b2: y = 16'hfe01;
			16'hf6b3: y = 16'hfe01;
			16'hf6b4: y = 16'hfe01;
			16'hf6b5: y = 16'hfe01;
			16'hf6b6: y = 16'hfe01;
			16'hf6b7: y = 16'hfe01;
			16'hf6b8: y = 16'hfe01;
			16'hf6b9: y = 16'hfe01;
			16'hf6ba: y = 16'hfe01;
			16'hf6bb: y = 16'hfe01;
			16'hf6bc: y = 16'hfe01;
			16'hf6bd: y = 16'hfe01;
			16'hf6be: y = 16'hfe01;
			16'hf6bf: y = 16'hfe01;
			16'hf6c0: y = 16'hfe01;
			16'hf6c1: y = 16'hfe01;
			16'hf6c2: y = 16'hfe01;
			16'hf6c3: y = 16'hfe01;
			16'hf6c4: y = 16'hfe01;
			16'hf6c5: y = 16'hfe01;
			16'hf6c6: y = 16'hfe01;
			16'hf6c7: y = 16'hfe01;
			16'hf6c8: y = 16'hfe01;
			16'hf6c9: y = 16'hfe01;
			16'hf6ca: y = 16'hfe01;
			16'hf6cb: y = 16'hfe01;
			16'hf6cc: y = 16'hfe01;
			16'hf6cd: y = 16'hfe01;
			16'hf6ce: y = 16'hfe01;
			16'hf6cf: y = 16'hfe01;
			16'hf6d0: y = 16'hfe01;
			16'hf6d1: y = 16'hfe01;
			16'hf6d2: y = 16'hfe01;
			16'hf6d3: y = 16'hfe01;
			16'hf6d4: y = 16'hfe01;
			16'hf6d5: y = 16'hfe01;
			16'hf6d6: y = 16'hfe01;
			16'hf6d7: y = 16'hfe01;
			16'hf6d8: y = 16'hfe01;
			16'hf6d9: y = 16'hfe01;
			16'hf6da: y = 16'hfe01;
			16'hf6db: y = 16'hfe01;
			16'hf6dc: y = 16'hfe01;
			16'hf6dd: y = 16'hfe01;
			16'hf6de: y = 16'hfe01;
			16'hf6df: y = 16'hfe01;
			16'hf6e0: y = 16'hfe01;
			16'hf6e1: y = 16'hfe01;
			16'hf6e2: y = 16'hfe01;
			16'hf6e3: y = 16'hfe01;
			16'hf6e4: y = 16'hfe01;
			16'hf6e5: y = 16'hfe01;
			16'hf6e6: y = 16'hfe01;
			16'hf6e7: y = 16'hfe01;
			16'hf6e8: y = 16'hfe01;
			16'hf6e9: y = 16'hfe01;
			16'hf6ea: y = 16'hfe01;
			16'hf6eb: y = 16'hfe01;
			16'hf6ec: y = 16'hfe01;
			16'hf6ed: y = 16'hfe01;
			16'hf6ee: y = 16'hfe01;
			16'hf6ef: y = 16'hfe01;
			16'hf6f0: y = 16'hfe01;
			16'hf6f1: y = 16'hfe01;
			16'hf6f2: y = 16'hfe01;
			16'hf6f3: y = 16'hfe01;
			16'hf6f4: y = 16'hfe01;
			16'hf6f5: y = 16'hfe01;
			16'hf6f6: y = 16'hfe01;
			16'hf6f7: y = 16'hfe01;
			16'hf6f8: y = 16'hfe01;
			16'hf6f9: y = 16'hfe01;
			16'hf6fa: y = 16'hfe01;
			16'hf6fb: y = 16'hfe01;
			16'hf6fc: y = 16'hfe01;
			16'hf6fd: y = 16'hfe01;
			16'hf6fe: y = 16'hfe01;
			16'hf6ff: y = 16'hfe01;
			16'hf700: y = 16'hfe01;
			16'hf701: y = 16'hfe01;
			16'hf702: y = 16'hfe01;
			16'hf703: y = 16'hfe01;
			16'hf704: y = 16'hfe01;
			16'hf705: y = 16'hfe01;
			16'hf706: y = 16'hfe01;
			16'hf707: y = 16'hfe01;
			16'hf708: y = 16'hfe01;
			16'hf709: y = 16'hfe01;
			16'hf70a: y = 16'hfe01;
			16'hf70b: y = 16'hfe01;
			16'hf70c: y = 16'hfe01;
			16'hf70d: y = 16'hfe01;
			16'hf70e: y = 16'hfe01;
			16'hf70f: y = 16'hfe01;
			16'hf710: y = 16'hfe01;
			16'hf711: y = 16'hfe01;
			16'hf712: y = 16'hfe01;
			16'hf713: y = 16'hfe01;
			16'hf714: y = 16'hfe01;
			16'hf715: y = 16'hfe01;
			16'hf716: y = 16'hfe01;
			16'hf717: y = 16'hfe01;
			16'hf718: y = 16'hfe01;
			16'hf719: y = 16'hfe01;
			16'hf71a: y = 16'hfe01;
			16'hf71b: y = 16'hfe01;
			16'hf71c: y = 16'hfe01;
			16'hf71d: y = 16'hfe01;
			16'hf71e: y = 16'hfe01;
			16'hf71f: y = 16'hfe01;
			16'hf720: y = 16'hfe01;
			16'hf721: y = 16'hfe01;
			16'hf722: y = 16'hfe01;
			16'hf723: y = 16'hfe01;
			16'hf724: y = 16'hfe01;
			16'hf725: y = 16'hfe01;
			16'hf726: y = 16'hfe01;
			16'hf727: y = 16'hfe01;
			16'hf728: y = 16'hfe01;
			16'hf729: y = 16'hfe01;
			16'hf72a: y = 16'hfe01;
			16'hf72b: y = 16'hfe01;
			16'hf72c: y = 16'hfe01;
			16'hf72d: y = 16'hfe01;
			16'hf72e: y = 16'hfe01;
			16'hf72f: y = 16'hfe01;
			16'hf730: y = 16'hfe01;
			16'hf731: y = 16'hfe01;
			16'hf732: y = 16'hfe01;
			16'hf733: y = 16'hfe01;
			16'hf734: y = 16'hfe01;
			16'hf735: y = 16'hfe01;
			16'hf736: y = 16'hfe01;
			16'hf737: y = 16'hfe01;
			16'hf738: y = 16'hfe01;
			16'hf739: y = 16'hfe01;
			16'hf73a: y = 16'hfe01;
			16'hf73b: y = 16'hfe01;
			16'hf73c: y = 16'hfe01;
			16'hf73d: y = 16'hfe01;
			16'hf73e: y = 16'hfe01;
			16'hf73f: y = 16'hfe01;
			16'hf740: y = 16'hfe01;
			16'hf741: y = 16'hfe01;
			16'hf742: y = 16'hfe01;
			16'hf743: y = 16'hfe01;
			16'hf744: y = 16'hfe01;
			16'hf745: y = 16'hfe01;
			16'hf746: y = 16'hfe01;
			16'hf747: y = 16'hfe01;
			16'hf748: y = 16'hfe01;
			16'hf749: y = 16'hfe01;
			16'hf74a: y = 16'hfe01;
			16'hf74b: y = 16'hfe01;
			16'hf74c: y = 16'hfe01;
			16'hf74d: y = 16'hfe01;
			16'hf74e: y = 16'hfe01;
			16'hf74f: y = 16'hfe01;
			16'hf750: y = 16'hfe01;
			16'hf751: y = 16'hfe01;
			16'hf752: y = 16'hfe01;
			16'hf753: y = 16'hfe01;
			16'hf754: y = 16'hfe01;
			16'hf755: y = 16'hfe01;
			16'hf756: y = 16'hfe01;
			16'hf757: y = 16'hfe01;
			16'hf758: y = 16'hfe01;
			16'hf759: y = 16'hfe01;
			16'hf75a: y = 16'hfe01;
			16'hf75b: y = 16'hfe01;
			16'hf75c: y = 16'hfe01;
			16'hf75d: y = 16'hfe01;
			16'hf75e: y = 16'hfe01;
			16'hf75f: y = 16'hfe01;
			16'hf760: y = 16'hfe01;
			16'hf761: y = 16'hfe01;
			16'hf762: y = 16'hfe01;
			16'hf763: y = 16'hfe01;
			16'hf764: y = 16'hfe01;
			16'hf765: y = 16'hfe01;
			16'hf766: y = 16'hfe01;
			16'hf767: y = 16'hfe01;
			16'hf768: y = 16'hfe01;
			16'hf769: y = 16'hfe01;
			16'hf76a: y = 16'hfe01;
			16'hf76b: y = 16'hfe01;
			16'hf76c: y = 16'hfe01;
			16'hf76d: y = 16'hfe01;
			16'hf76e: y = 16'hfe01;
			16'hf76f: y = 16'hfe01;
			16'hf770: y = 16'hfe01;
			16'hf771: y = 16'hfe01;
			16'hf772: y = 16'hfe01;
			16'hf773: y = 16'hfe01;
			16'hf774: y = 16'hfe01;
			16'hf775: y = 16'hfe01;
			16'hf776: y = 16'hfe01;
			16'hf777: y = 16'hfe01;
			16'hf778: y = 16'hfe01;
			16'hf779: y = 16'hfe01;
			16'hf77a: y = 16'hfe01;
			16'hf77b: y = 16'hfe01;
			16'hf77c: y = 16'hfe01;
			16'hf77d: y = 16'hfe01;
			16'hf77e: y = 16'hfe01;
			16'hf77f: y = 16'hfe01;
			16'hf780: y = 16'hfe01;
			16'hf781: y = 16'hfe01;
			16'hf782: y = 16'hfe01;
			16'hf783: y = 16'hfe01;
			16'hf784: y = 16'hfe01;
			16'hf785: y = 16'hfe01;
			16'hf786: y = 16'hfe01;
			16'hf787: y = 16'hfe01;
			16'hf788: y = 16'hfe01;
			16'hf789: y = 16'hfe01;
			16'hf78a: y = 16'hfe01;
			16'hf78b: y = 16'hfe01;
			16'hf78c: y = 16'hfe01;
			16'hf78d: y = 16'hfe01;
			16'hf78e: y = 16'hfe01;
			16'hf78f: y = 16'hfe01;
			16'hf790: y = 16'hfe01;
			16'hf791: y = 16'hfe01;
			16'hf792: y = 16'hfe01;
			16'hf793: y = 16'hfe01;
			16'hf794: y = 16'hfe01;
			16'hf795: y = 16'hfe01;
			16'hf796: y = 16'hfe01;
			16'hf797: y = 16'hfe01;
			16'hf798: y = 16'hfe01;
			16'hf799: y = 16'hfe01;
			16'hf79a: y = 16'hfe01;
			16'hf79b: y = 16'hfe01;
			16'hf79c: y = 16'hfe01;
			16'hf79d: y = 16'hfe01;
			16'hf79e: y = 16'hfe01;
			16'hf79f: y = 16'hfe01;
			16'hf7a0: y = 16'hfe01;
			16'hf7a1: y = 16'hfe01;
			16'hf7a2: y = 16'hfe01;
			16'hf7a3: y = 16'hfe01;
			16'hf7a4: y = 16'hfe01;
			16'hf7a5: y = 16'hfe01;
			16'hf7a6: y = 16'hfe01;
			16'hf7a7: y = 16'hfe01;
			16'hf7a8: y = 16'hfe01;
			16'hf7a9: y = 16'hfe01;
			16'hf7aa: y = 16'hfe01;
			16'hf7ab: y = 16'hfe01;
			16'hf7ac: y = 16'hfe01;
			16'hf7ad: y = 16'hfe01;
			16'hf7ae: y = 16'hfe01;
			16'hf7af: y = 16'hfe01;
			16'hf7b0: y = 16'hfe01;
			16'hf7b1: y = 16'hfe01;
			16'hf7b2: y = 16'hfe01;
			16'hf7b3: y = 16'hfe01;
			16'hf7b4: y = 16'hfe01;
			16'hf7b5: y = 16'hfe01;
			16'hf7b6: y = 16'hfe01;
			16'hf7b7: y = 16'hfe01;
			16'hf7b8: y = 16'hfe01;
			16'hf7b9: y = 16'hfe01;
			16'hf7ba: y = 16'hfe01;
			16'hf7bb: y = 16'hfe01;
			16'hf7bc: y = 16'hfe01;
			16'hf7bd: y = 16'hfe01;
			16'hf7be: y = 16'hfe01;
			16'hf7bf: y = 16'hfe01;
			16'hf7c0: y = 16'hfe01;
			16'hf7c1: y = 16'hfe01;
			16'hf7c2: y = 16'hfe01;
			16'hf7c3: y = 16'hfe01;
			16'hf7c4: y = 16'hfe01;
			16'hf7c5: y = 16'hfe01;
			16'hf7c6: y = 16'hfe01;
			16'hf7c7: y = 16'hfe01;
			16'hf7c8: y = 16'hfe01;
			16'hf7c9: y = 16'hfe01;
			16'hf7ca: y = 16'hfe01;
			16'hf7cb: y = 16'hfe01;
			16'hf7cc: y = 16'hfe01;
			16'hf7cd: y = 16'hfe01;
			16'hf7ce: y = 16'hfe01;
			16'hf7cf: y = 16'hfe01;
			16'hf7d0: y = 16'hfe01;
			16'hf7d1: y = 16'hfe01;
			16'hf7d2: y = 16'hfe01;
			16'hf7d3: y = 16'hfe01;
			16'hf7d4: y = 16'hfe01;
			16'hf7d5: y = 16'hfe01;
			16'hf7d6: y = 16'hfe01;
			16'hf7d7: y = 16'hfe01;
			16'hf7d8: y = 16'hfe01;
			16'hf7d9: y = 16'hfe01;
			16'hf7da: y = 16'hfe01;
			16'hf7db: y = 16'hfe01;
			16'hf7dc: y = 16'hfe01;
			16'hf7dd: y = 16'hfe01;
			16'hf7de: y = 16'hfe01;
			16'hf7df: y = 16'hfe01;
			16'hf7e0: y = 16'hfe01;
			16'hf7e1: y = 16'hfe01;
			16'hf7e2: y = 16'hfe01;
			16'hf7e3: y = 16'hfe01;
			16'hf7e4: y = 16'hfe01;
			16'hf7e5: y = 16'hfe01;
			16'hf7e6: y = 16'hfe01;
			16'hf7e7: y = 16'hfe01;
			16'hf7e8: y = 16'hfe01;
			16'hf7e9: y = 16'hfe01;
			16'hf7ea: y = 16'hfe01;
			16'hf7eb: y = 16'hfe01;
			16'hf7ec: y = 16'hfe01;
			16'hf7ed: y = 16'hfe01;
			16'hf7ee: y = 16'hfe01;
			16'hf7ef: y = 16'hfe01;
			16'hf7f0: y = 16'hfe01;
			16'hf7f1: y = 16'hfe01;
			16'hf7f2: y = 16'hfe01;
			16'hf7f3: y = 16'hfe01;
			16'hf7f4: y = 16'hfe01;
			16'hf7f5: y = 16'hfe01;
			16'hf7f6: y = 16'hfe01;
			16'hf7f7: y = 16'hfe01;
			16'hf7f8: y = 16'hfe01;
			16'hf7f9: y = 16'hfe01;
			16'hf7fa: y = 16'hfe01;
			16'hf7fb: y = 16'hfe01;
			16'hf7fc: y = 16'hfe01;
			16'hf7fd: y = 16'hfe01;
			16'hf7fe: y = 16'hfe01;
			16'hf7ff: y = 16'hfe01;
			16'hf800: y = 16'hfe01;
			16'hf801: y = 16'hfe01;
			16'hf802: y = 16'hfe01;
			16'hf803: y = 16'hfe01;
			16'hf804: y = 16'hfe01;
			16'hf805: y = 16'hfe01;
			16'hf806: y = 16'hfe01;
			16'hf807: y = 16'hfe01;
			16'hf808: y = 16'hfe01;
			16'hf809: y = 16'hfe01;
			16'hf80a: y = 16'hfe01;
			16'hf80b: y = 16'hfe01;
			16'hf80c: y = 16'hfe01;
			16'hf80d: y = 16'hfe01;
			16'hf80e: y = 16'hfe01;
			16'hf80f: y = 16'hfe01;
			16'hf810: y = 16'hfe01;
			16'hf811: y = 16'hfe01;
			16'hf812: y = 16'hfe01;
			16'hf813: y = 16'hfe01;
			16'hf814: y = 16'hfe01;
			16'hf815: y = 16'hfe01;
			16'hf816: y = 16'hfe01;
			16'hf817: y = 16'hfe01;
			16'hf818: y = 16'hfe01;
			16'hf819: y = 16'hfe01;
			16'hf81a: y = 16'hfe01;
			16'hf81b: y = 16'hfe01;
			16'hf81c: y = 16'hfe01;
			16'hf81d: y = 16'hfe01;
			16'hf81e: y = 16'hfe01;
			16'hf81f: y = 16'hfe01;
			16'hf820: y = 16'hfe01;
			16'hf821: y = 16'hfe01;
			16'hf822: y = 16'hfe01;
			16'hf823: y = 16'hfe01;
			16'hf824: y = 16'hfe01;
			16'hf825: y = 16'hfe01;
			16'hf826: y = 16'hfe01;
			16'hf827: y = 16'hfe01;
			16'hf828: y = 16'hfe01;
			16'hf829: y = 16'hfe01;
			16'hf82a: y = 16'hfe01;
			16'hf82b: y = 16'hfe01;
			16'hf82c: y = 16'hfe01;
			16'hf82d: y = 16'hfe01;
			16'hf82e: y = 16'hfe01;
			16'hf82f: y = 16'hfe01;
			16'hf830: y = 16'hfe01;
			16'hf831: y = 16'hfe01;
			16'hf832: y = 16'hfe01;
			16'hf833: y = 16'hfe01;
			16'hf834: y = 16'hfe01;
			16'hf835: y = 16'hfe01;
			16'hf836: y = 16'hfe01;
			16'hf837: y = 16'hfe01;
			16'hf838: y = 16'hfe01;
			16'hf839: y = 16'hfe01;
			16'hf83a: y = 16'hfe01;
			16'hf83b: y = 16'hfe01;
			16'hf83c: y = 16'hfe01;
			16'hf83d: y = 16'hfe01;
			16'hf83e: y = 16'hfe01;
			16'hf83f: y = 16'hfe01;
			16'hf840: y = 16'hfe01;
			16'hf841: y = 16'hfe01;
			16'hf842: y = 16'hfe01;
			16'hf843: y = 16'hfe01;
			16'hf844: y = 16'hfe01;
			16'hf845: y = 16'hfe01;
			16'hf846: y = 16'hfe01;
			16'hf847: y = 16'hfe01;
			16'hf848: y = 16'hfe01;
			16'hf849: y = 16'hfe01;
			16'hf84a: y = 16'hfe01;
			16'hf84b: y = 16'hfe01;
			16'hf84c: y = 16'hfe01;
			16'hf84d: y = 16'hfe01;
			16'hf84e: y = 16'hfe01;
			16'hf84f: y = 16'hfe01;
			16'hf850: y = 16'hfe01;
			16'hf851: y = 16'hfe01;
			16'hf852: y = 16'hfe01;
			16'hf853: y = 16'hfe01;
			16'hf854: y = 16'hfe01;
			16'hf855: y = 16'hfe01;
			16'hf856: y = 16'hfe01;
			16'hf857: y = 16'hfe01;
			16'hf858: y = 16'hfe01;
			16'hf859: y = 16'hfe01;
			16'hf85a: y = 16'hfe01;
			16'hf85b: y = 16'hfe01;
			16'hf85c: y = 16'hfe01;
			16'hf85d: y = 16'hfe01;
			16'hf85e: y = 16'hfe01;
			16'hf85f: y = 16'hfe01;
			16'hf860: y = 16'hfe01;
			16'hf861: y = 16'hfe01;
			16'hf862: y = 16'hfe01;
			16'hf863: y = 16'hfe01;
			16'hf864: y = 16'hfe01;
			16'hf865: y = 16'hfe01;
			16'hf866: y = 16'hfe01;
			16'hf867: y = 16'hfe01;
			16'hf868: y = 16'hfe01;
			16'hf869: y = 16'hfe01;
			16'hf86a: y = 16'hfe01;
			16'hf86b: y = 16'hfe01;
			16'hf86c: y = 16'hfe01;
			16'hf86d: y = 16'hfe01;
			16'hf86e: y = 16'hfe01;
			16'hf86f: y = 16'hfe01;
			16'hf870: y = 16'hfe01;
			16'hf871: y = 16'hfe01;
			16'hf872: y = 16'hfe01;
			16'hf873: y = 16'hfe01;
			16'hf874: y = 16'hfe01;
			16'hf875: y = 16'hfe01;
			16'hf876: y = 16'hfe01;
			16'hf877: y = 16'hfe01;
			16'hf878: y = 16'hfe01;
			16'hf879: y = 16'hfe01;
			16'hf87a: y = 16'hfe01;
			16'hf87b: y = 16'hfe01;
			16'hf87c: y = 16'hfe01;
			16'hf87d: y = 16'hfe01;
			16'hf87e: y = 16'hfe01;
			16'hf87f: y = 16'hfe01;
			16'hf880: y = 16'hfe01;
			16'hf881: y = 16'hfe01;
			16'hf882: y = 16'hfe01;
			16'hf883: y = 16'hfe01;
			16'hf884: y = 16'hfe01;
			16'hf885: y = 16'hfe01;
			16'hf886: y = 16'hfe01;
			16'hf887: y = 16'hfe01;
			16'hf888: y = 16'hfe01;
			16'hf889: y = 16'hfe01;
			16'hf88a: y = 16'hfe01;
			16'hf88b: y = 16'hfe01;
			16'hf88c: y = 16'hfe01;
			16'hf88d: y = 16'hfe01;
			16'hf88e: y = 16'hfe01;
			16'hf88f: y = 16'hfe01;
			16'hf890: y = 16'hfe01;
			16'hf891: y = 16'hfe01;
			16'hf892: y = 16'hfe01;
			16'hf893: y = 16'hfe01;
			16'hf894: y = 16'hfe01;
			16'hf895: y = 16'hfe01;
			16'hf896: y = 16'hfe01;
			16'hf897: y = 16'hfe01;
			16'hf898: y = 16'hfe01;
			16'hf899: y = 16'hfe01;
			16'hf89a: y = 16'hfe01;
			16'hf89b: y = 16'hfe01;
			16'hf89c: y = 16'hfe01;
			16'hf89d: y = 16'hfe01;
			16'hf89e: y = 16'hfe01;
			16'hf89f: y = 16'hfe01;
			16'hf8a0: y = 16'hfe01;
			16'hf8a1: y = 16'hfe01;
			16'hf8a2: y = 16'hfe01;
			16'hf8a3: y = 16'hfe01;
			16'hf8a4: y = 16'hfe01;
			16'hf8a5: y = 16'hfe01;
			16'hf8a6: y = 16'hfe01;
			16'hf8a7: y = 16'hfe01;
			16'hf8a8: y = 16'hfe01;
			16'hf8a9: y = 16'hfe01;
			16'hf8aa: y = 16'hfe01;
			16'hf8ab: y = 16'hfe01;
			16'hf8ac: y = 16'hfe01;
			16'hf8ad: y = 16'hfe01;
			16'hf8ae: y = 16'hfe01;
			16'hf8af: y = 16'hfe01;
			16'hf8b0: y = 16'hfe01;
			16'hf8b1: y = 16'hfe01;
			16'hf8b2: y = 16'hfe01;
			16'hf8b3: y = 16'hfe01;
			16'hf8b4: y = 16'hfe01;
			16'hf8b5: y = 16'hfe01;
			16'hf8b6: y = 16'hfe01;
			16'hf8b7: y = 16'hfe01;
			16'hf8b8: y = 16'hfe01;
			16'hf8b9: y = 16'hfe01;
			16'hf8ba: y = 16'hfe01;
			16'hf8bb: y = 16'hfe01;
			16'hf8bc: y = 16'hfe01;
			16'hf8bd: y = 16'hfe01;
			16'hf8be: y = 16'hfe01;
			16'hf8bf: y = 16'hfe01;
			16'hf8c0: y = 16'hfe01;
			16'hf8c1: y = 16'hfe01;
			16'hf8c2: y = 16'hfe01;
			16'hf8c3: y = 16'hfe01;
			16'hf8c4: y = 16'hfe01;
			16'hf8c5: y = 16'hfe01;
			16'hf8c6: y = 16'hfe01;
			16'hf8c7: y = 16'hfe01;
			16'hf8c8: y = 16'hfe01;
			16'hf8c9: y = 16'hfe01;
			16'hf8ca: y = 16'hfe01;
			16'hf8cb: y = 16'hfe01;
			16'hf8cc: y = 16'hfe01;
			16'hf8cd: y = 16'hfe01;
			16'hf8ce: y = 16'hfe01;
			16'hf8cf: y = 16'hfe01;
			16'hf8d0: y = 16'hfe01;
			16'hf8d1: y = 16'hfe01;
			16'hf8d2: y = 16'hfe01;
			16'hf8d3: y = 16'hfe01;
			16'hf8d4: y = 16'hfe01;
			16'hf8d5: y = 16'hfe01;
			16'hf8d6: y = 16'hfe01;
			16'hf8d7: y = 16'hfe01;
			16'hf8d8: y = 16'hfe01;
			16'hf8d9: y = 16'hfe01;
			16'hf8da: y = 16'hfe01;
			16'hf8db: y = 16'hfe01;
			16'hf8dc: y = 16'hfe01;
			16'hf8dd: y = 16'hfe01;
			16'hf8de: y = 16'hfe01;
			16'hf8df: y = 16'hfe01;
			16'hf8e0: y = 16'hfe01;
			16'hf8e1: y = 16'hfe01;
			16'hf8e2: y = 16'hfe01;
			16'hf8e3: y = 16'hfe01;
			16'hf8e4: y = 16'hfe01;
			16'hf8e5: y = 16'hfe01;
			16'hf8e6: y = 16'hfe01;
			16'hf8e7: y = 16'hfe01;
			16'hf8e8: y = 16'hfe01;
			16'hf8e9: y = 16'hfe01;
			16'hf8ea: y = 16'hfe01;
			16'hf8eb: y = 16'hfe01;
			16'hf8ec: y = 16'hfe01;
			16'hf8ed: y = 16'hfe01;
			16'hf8ee: y = 16'hfe01;
			16'hf8ef: y = 16'hfe01;
			16'hf8f0: y = 16'hfe01;
			16'hf8f1: y = 16'hfe01;
			16'hf8f2: y = 16'hfe01;
			16'hf8f3: y = 16'hfe01;
			16'hf8f4: y = 16'hfe01;
			16'hf8f5: y = 16'hfe01;
			16'hf8f6: y = 16'hfe01;
			16'hf8f7: y = 16'hfe01;
			16'hf8f8: y = 16'hfe01;
			16'hf8f9: y = 16'hfe01;
			16'hf8fa: y = 16'hfe01;
			16'hf8fb: y = 16'hfe01;
			16'hf8fc: y = 16'hfe01;
			16'hf8fd: y = 16'hfe01;
			16'hf8fe: y = 16'hfe01;
			16'hf8ff: y = 16'hfe01;
			16'hf900: y = 16'hfe01;
			16'hf901: y = 16'hfe01;
			16'hf902: y = 16'hfe01;
			16'hf903: y = 16'hfe01;
			16'hf904: y = 16'hfe01;
			16'hf905: y = 16'hfe01;
			16'hf906: y = 16'hfe01;
			16'hf907: y = 16'hfe01;
			16'hf908: y = 16'hfe01;
			16'hf909: y = 16'hfe01;
			16'hf90a: y = 16'hfe01;
			16'hf90b: y = 16'hfe01;
			16'hf90c: y = 16'hfe01;
			16'hf90d: y = 16'hfe01;
			16'hf90e: y = 16'hfe01;
			16'hf90f: y = 16'hfe01;
			16'hf910: y = 16'hfe01;
			16'hf911: y = 16'hfe01;
			16'hf912: y = 16'hfe02;
			16'hf913: y = 16'hfe02;
			16'hf914: y = 16'hfe02;
			16'hf915: y = 16'hfe02;
			16'hf916: y = 16'hfe02;
			16'hf917: y = 16'hfe02;
			16'hf918: y = 16'hfe02;
			16'hf919: y = 16'hfe02;
			16'hf91a: y = 16'hfe02;
			16'hf91b: y = 16'hfe02;
			16'hf91c: y = 16'hfe02;
			16'hf91d: y = 16'hfe02;
			16'hf91e: y = 16'hfe02;
			16'hf91f: y = 16'hfe02;
			16'hf920: y = 16'hfe02;
			16'hf921: y = 16'hfe02;
			16'hf922: y = 16'hfe02;
			16'hf923: y = 16'hfe02;
			16'hf924: y = 16'hfe02;
			16'hf925: y = 16'hfe02;
			16'hf926: y = 16'hfe02;
			16'hf927: y = 16'hfe02;
			16'hf928: y = 16'hfe02;
			16'hf929: y = 16'hfe02;
			16'hf92a: y = 16'hfe02;
			16'hf92b: y = 16'hfe02;
			16'hf92c: y = 16'hfe02;
			16'hf92d: y = 16'hfe02;
			16'hf92e: y = 16'hfe02;
			16'hf92f: y = 16'hfe02;
			16'hf930: y = 16'hfe02;
			16'hf931: y = 16'hfe02;
			16'hf932: y = 16'hfe02;
			16'hf933: y = 16'hfe02;
			16'hf934: y = 16'hfe02;
			16'hf935: y = 16'hfe02;
			16'hf936: y = 16'hfe02;
			16'hf937: y = 16'hfe02;
			16'hf938: y = 16'hfe02;
			16'hf939: y = 16'hfe02;
			16'hf93a: y = 16'hfe02;
			16'hf93b: y = 16'hfe02;
			16'hf93c: y = 16'hfe02;
			16'hf93d: y = 16'hfe02;
			16'hf93e: y = 16'hfe02;
			16'hf93f: y = 16'hfe02;
			16'hf940: y = 16'hfe02;
			16'hf941: y = 16'hfe02;
			16'hf942: y = 16'hfe02;
			16'hf943: y = 16'hfe02;
			16'hf944: y = 16'hfe02;
			16'hf945: y = 16'hfe02;
			16'hf946: y = 16'hfe02;
			16'hf947: y = 16'hfe02;
			16'hf948: y = 16'hfe02;
			16'hf949: y = 16'hfe02;
			16'hf94a: y = 16'hfe02;
			16'hf94b: y = 16'hfe02;
			16'hf94c: y = 16'hfe02;
			16'hf94d: y = 16'hfe02;
			16'hf94e: y = 16'hfe02;
			16'hf94f: y = 16'hfe02;
			16'hf950: y = 16'hfe02;
			16'hf951: y = 16'hfe02;
			16'hf952: y = 16'hfe02;
			16'hf953: y = 16'hfe02;
			16'hf954: y = 16'hfe02;
			16'hf955: y = 16'hfe02;
			16'hf956: y = 16'hfe02;
			16'hf957: y = 16'hfe02;
			16'hf958: y = 16'hfe02;
			16'hf959: y = 16'hfe02;
			16'hf95a: y = 16'hfe02;
			16'hf95b: y = 16'hfe02;
			16'hf95c: y = 16'hfe02;
			16'hf95d: y = 16'hfe02;
			16'hf95e: y = 16'hfe02;
			16'hf95f: y = 16'hfe02;
			16'hf960: y = 16'hfe02;
			16'hf961: y = 16'hfe02;
			16'hf962: y = 16'hfe02;
			16'hf963: y = 16'hfe02;
			16'hf964: y = 16'hfe02;
			16'hf965: y = 16'hfe02;
			16'hf966: y = 16'hfe02;
			16'hf967: y = 16'hfe02;
			16'hf968: y = 16'hfe02;
			16'hf969: y = 16'hfe02;
			16'hf96a: y = 16'hfe02;
			16'hf96b: y = 16'hfe02;
			16'hf96c: y = 16'hfe02;
			16'hf96d: y = 16'hfe02;
			16'hf96e: y = 16'hfe02;
			16'hf96f: y = 16'hfe02;
			16'hf970: y = 16'hfe02;
			16'hf971: y = 16'hfe02;
			16'hf972: y = 16'hfe02;
			16'hf973: y = 16'hfe02;
			16'hf974: y = 16'hfe02;
			16'hf975: y = 16'hfe02;
			16'hf976: y = 16'hfe02;
			16'hf977: y = 16'hfe02;
			16'hf978: y = 16'hfe02;
			16'hf979: y = 16'hfe02;
			16'hf97a: y = 16'hfe02;
			16'hf97b: y = 16'hfe02;
			16'hf97c: y = 16'hfe02;
			16'hf97d: y = 16'hfe02;
			16'hf97e: y = 16'hfe02;
			16'hf97f: y = 16'hfe02;
			16'hf980: y = 16'hfe02;
			16'hf981: y = 16'hfe02;
			16'hf982: y = 16'hfe02;
			16'hf983: y = 16'hfe02;
			16'hf984: y = 16'hfe02;
			16'hf985: y = 16'hfe02;
			16'hf986: y = 16'hfe02;
			16'hf987: y = 16'hfe02;
			16'hf988: y = 16'hfe02;
			16'hf989: y = 16'hfe02;
			16'hf98a: y = 16'hfe02;
			16'hf98b: y = 16'hfe02;
			16'hf98c: y = 16'hfe02;
			16'hf98d: y = 16'hfe02;
			16'hf98e: y = 16'hfe02;
			16'hf98f: y = 16'hfe02;
			16'hf990: y = 16'hfe02;
			16'hf991: y = 16'hfe02;
			16'hf992: y = 16'hfe02;
			16'hf993: y = 16'hfe02;
			16'hf994: y = 16'hfe02;
			16'hf995: y = 16'hfe02;
			16'hf996: y = 16'hfe02;
			16'hf997: y = 16'hfe02;
			16'hf998: y = 16'hfe02;
			16'hf999: y = 16'hfe02;
			16'hf99a: y = 16'hfe02;
			16'hf99b: y = 16'hfe02;
			16'hf99c: y = 16'hfe02;
			16'hf99d: y = 16'hfe02;
			16'hf99e: y = 16'hfe02;
			16'hf99f: y = 16'hfe02;
			16'hf9a0: y = 16'hfe02;
			16'hf9a1: y = 16'hfe02;
			16'hf9a2: y = 16'hfe02;
			16'hf9a3: y = 16'hfe02;
			16'hf9a4: y = 16'hfe02;
			16'hf9a5: y = 16'hfe02;
			16'hf9a6: y = 16'hfe02;
			16'hf9a7: y = 16'hfe02;
			16'hf9a8: y = 16'hfe02;
			16'hf9a9: y = 16'hfe02;
			16'hf9aa: y = 16'hfe02;
			16'hf9ab: y = 16'hfe02;
			16'hf9ac: y = 16'hfe02;
			16'hf9ad: y = 16'hfe02;
			16'hf9ae: y = 16'hfe02;
			16'hf9af: y = 16'hfe02;
			16'hf9b0: y = 16'hfe02;
			16'hf9b1: y = 16'hfe02;
			16'hf9b2: y = 16'hfe02;
			16'hf9b3: y = 16'hfe02;
			16'hf9b4: y = 16'hfe02;
			16'hf9b5: y = 16'hfe02;
			16'hf9b6: y = 16'hfe02;
			16'hf9b7: y = 16'hfe02;
			16'hf9b8: y = 16'hfe02;
			16'hf9b9: y = 16'hfe02;
			16'hf9ba: y = 16'hfe02;
			16'hf9bb: y = 16'hfe02;
			16'hf9bc: y = 16'hfe02;
			16'hf9bd: y = 16'hfe02;
			16'hf9be: y = 16'hfe02;
			16'hf9bf: y = 16'hfe02;
			16'hf9c0: y = 16'hfe02;
			16'hf9c1: y = 16'hfe02;
			16'hf9c2: y = 16'hfe02;
			16'hf9c3: y = 16'hfe02;
			16'hf9c4: y = 16'hfe03;
			16'hf9c5: y = 16'hfe03;
			16'hf9c6: y = 16'hfe03;
			16'hf9c7: y = 16'hfe03;
			16'hf9c8: y = 16'hfe03;
			16'hf9c9: y = 16'hfe03;
			16'hf9ca: y = 16'hfe03;
			16'hf9cb: y = 16'hfe03;
			16'hf9cc: y = 16'hfe03;
			16'hf9cd: y = 16'hfe03;
			16'hf9ce: y = 16'hfe03;
			16'hf9cf: y = 16'hfe03;
			16'hf9d0: y = 16'hfe03;
			16'hf9d1: y = 16'hfe03;
			16'hf9d2: y = 16'hfe03;
			16'hf9d3: y = 16'hfe03;
			16'hf9d4: y = 16'hfe03;
			16'hf9d5: y = 16'hfe03;
			16'hf9d6: y = 16'hfe03;
			16'hf9d7: y = 16'hfe03;
			16'hf9d8: y = 16'hfe03;
			16'hf9d9: y = 16'hfe03;
			16'hf9da: y = 16'hfe03;
			16'hf9db: y = 16'hfe03;
			16'hf9dc: y = 16'hfe03;
			16'hf9dd: y = 16'hfe03;
			16'hf9de: y = 16'hfe03;
			16'hf9df: y = 16'hfe03;
			16'hf9e0: y = 16'hfe03;
			16'hf9e1: y = 16'hfe03;
			16'hf9e2: y = 16'hfe03;
			16'hf9e3: y = 16'hfe03;
			16'hf9e4: y = 16'hfe03;
			16'hf9e5: y = 16'hfe03;
			16'hf9e6: y = 16'hfe03;
			16'hf9e7: y = 16'hfe03;
			16'hf9e8: y = 16'hfe03;
			16'hf9e9: y = 16'hfe03;
			16'hf9ea: y = 16'hfe03;
			16'hf9eb: y = 16'hfe03;
			16'hf9ec: y = 16'hfe03;
			16'hf9ed: y = 16'hfe03;
			16'hf9ee: y = 16'hfe03;
			16'hf9ef: y = 16'hfe03;
			16'hf9f0: y = 16'hfe03;
			16'hf9f1: y = 16'hfe03;
			16'hf9f2: y = 16'hfe03;
			16'hf9f3: y = 16'hfe03;
			16'hf9f4: y = 16'hfe03;
			16'hf9f5: y = 16'hfe03;
			16'hf9f6: y = 16'hfe03;
			16'hf9f7: y = 16'hfe03;
			16'hf9f8: y = 16'hfe03;
			16'hf9f9: y = 16'hfe03;
			16'hf9fa: y = 16'hfe03;
			16'hf9fb: y = 16'hfe03;
			16'hf9fc: y = 16'hfe03;
			16'hf9fd: y = 16'hfe03;
			16'hf9fe: y = 16'hfe03;
			16'hf9ff: y = 16'hfe03;
			16'hfa00: y = 16'hfe03;
			16'hfa01: y = 16'hfe03;
			16'hfa02: y = 16'hfe03;
			16'hfa03: y = 16'hfe03;
			16'hfa04: y = 16'hfe03;
			16'hfa05: y = 16'hfe03;
			16'hfa06: y = 16'hfe03;
			16'hfa07: y = 16'hfe03;
			16'hfa08: y = 16'hfe03;
			16'hfa09: y = 16'hfe03;
			16'hfa0a: y = 16'hfe03;
			16'hfa0b: y = 16'hfe03;
			16'hfa0c: y = 16'hfe03;
			16'hfa0d: y = 16'hfe03;
			16'hfa0e: y = 16'hfe03;
			16'hfa0f: y = 16'hfe03;
			16'hfa10: y = 16'hfe03;
			16'hfa11: y = 16'hfe03;
			16'hfa12: y = 16'hfe03;
			16'hfa13: y = 16'hfe03;
			16'hfa14: y = 16'hfe03;
			16'hfa15: y = 16'hfe03;
			16'hfa16: y = 16'hfe03;
			16'hfa17: y = 16'hfe03;
			16'hfa18: y = 16'hfe03;
			16'hfa19: y = 16'hfe03;
			16'hfa1a: y = 16'hfe03;
			16'hfa1b: y = 16'hfe03;
			16'hfa1c: y = 16'hfe03;
			16'hfa1d: y = 16'hfe03;
			16'hfa1e: y = 16'hfe03;
			16'hfa1f: y = 16'hfe03;
			16'hfa20: y = 16'hfe03;
			16'hfa21: y = 16'hfe03;
			16'hfa22: y = 16'hfe03;
			16'hfa23: y = 16'hfe03;
			16'hfa24: y = 16'hfe03;
			16'hfa25: y = 16'hfe03;
			16'hfa26: y = 16'hfe03;
			16'hfa27: y = 16'hfe03;
			16'hfa28: y = 16'hfe03;
			16'hfa29: y = 16'hfe03;
			16'hfa2a: y = 16'hfe03;
			16'hfa2b: y = 16'hfe03;
			16'hfa2c: y = 16'hfe04;
			16'hfa2d: y = 16'hfe04;
			16'hfa2e: y = 16'hfe04;
			16'hfa2f: y = 16'hfe04;
			16'hfa30: y = 16'hfe04;
			16'hfa31: y = 16'hfe04;
			16'hfa32: y = 16'hfe04;
			16'hfa33: y = 16'hfe04;
			16'hfa34: y = 16'hfe04;
			16'hfa35: y = 16'hfe04;
			16'hfa36: y = 16'hfe04;
			16'hfa37: y = 16'hfe04;
			16'hfa38: y = 16'hfe04;
			16'hfa39: y = 16'hfe04;
			16'hfa3a: y = 16'hfe04;
			16'hfa3b: y = 16'hfe04;
			16'hfa3c: y = 16'hfe04;
			16'hfa3d: y = 16'hfe04;
			16'hfa3e: y = 16'hfe04;
			16'hfa3f: y = 16'hfe04;
			16'hfa40: y = 16'hfe04;
			16'hfa41: y = 16'hfe04;
			16'hfa42: y = 16'hfe04;
			16'hfa43: y = 16'hfe04;
			16'hfa44: y = 16'hfe04;
			16'hfa45: y = 16'hfe04;
			16'hfa46: y = 16'hfe04;
			16'hfa47: y = 16'hfe04;
			16'hfa48: y = 16'hfe04;
			16'hfa49: y = 16'hfe04;
			16'hfa4a: y = 16'hfe04;
			16'hfa4b: y = 16'hfe04;
			16'hfa4c: y = 16'hfe04;
			16'hfa4d: y = 16'hfe04;
			16'hfa4e: y = 16'hfe04;
			16'hfa4f: y = 16'hfe04;
			16'hfa50: y = 16'hfe04;
			16'hfa51: y = 16'hfe04;
			16'hfa52: y = 16'hfe04;
			16'hfa53: y = 16'hfe04;
			16'hfa54: y = 16'hfe04;
			16'hfa55: y = 16'hfe04;
			16'hfa56: y = 16'hfe04;
			16'hfa57: y = 16'hfe04;
			16'hfa58: y = 16'hfe04;
			16'hfa59: y = 16'hfe04;
			16'hfa5a: y = 16'hfe04;
			16'hfa5b: y = 16'hfe04;
			16'hfa5c: y = 16'hfe04;
			16'hfa5d: y = 16'hfe04;
			16'hfa5e: y = 16'hfe04;
			16'hfa5f: y = 16'hfe04;
			16'hfa60: y = 16'hfe04;
			16'hfa61: y = 16'hfe04;
			16'hfa62: y = 16'hfe04;
			16'hfa63: y = 16'hfe04;
			16'hfa64: y = 16'hfe04;
			16'hfa65: y = 16'hfe04;
			16'hfa66: y = 16'hfe04;
			16'hfa67: y = 16'hfe04;
			16'hfa68: y = 16'hfe04;
			16'hfa69: y = 16'hfe04;
			16'hfa6a: y = 16'hfe04;
			16'hfa6b: y = 16'hfe04;
			16'hfa6c: y = 16'hfe04;
			16'hfa6d: y = 16'hfe04;
			16'hfa6e: y = 16'hfe04;
			16'hfa6f: y = 16'hfe04;
			16'hfa70: y = 16'hfe04;
			16'hfa71: y = 16'hfe04;
			16'hfa72: y = 16'hfe04;
			16'hfa73: y = 16'hfe04;
			16'hfa74: y = 16'hfe04;
			16'hfa75: y = 16'hfe04;
			16'hfa76: y = 16'hfe05;
			16'hfa77: y = 16'hfe05;
			16'hfa78: y = 16'hfe05;
			16'hfa79: y = 16'hfe05;
			16'hfa7a: y = 16'hfe05;
			16'hfa7b: y = 16'hfe05;
			16'hfa7c: y = 16'hfe05;
			16'hfa7d: y = 16'hfe05;
			16'hfa7e: y = 16'hfe05;
			16'hfa7f: y = 16'hfe05;
			16'hfa80: y = 16'hfe05;
			16'hfa81: y = 16'hfe05;
			16'hfa82: y = 16'hfe05;
			16'hfa83: y = 16'hfe05;
			16'hfa84: y = 16'hfe05;
			16'hfa85: y = 16'hfe05;
			16'hfa86: y = 16'hfe05;
			16'hfa87: y = 16'hfe05;
			16'hfa88: y = 16'hfe05;
			16'hfa89: y = 16'hfe05;
			16'hfa8a: y = 16'hfe05;
			16'hfa8b: y = 16'hfe05;
			16'hfa8c: y = 16'hfe05;
			16'hfa8d: y = 16'hfe05;
			16'hfa8e: y = 16'hfe05;
			16'hfa8f: y = 16'hfe05;
			16'hfa90: y = 16'hfe05;
			16'hfa91: y = 16'hfe05;
			16'hfa92: y = 16'hfe05;
			16'hfa93: y = 16'hfe05;
			16'hfa94: y = 16'hfe05;
			16'hfa95: y = 16'hfe05;
			16'hfa96: y = 16'hfe05;
			16'hfa97: y = 16'hfe05;
			16'hfa98: y = 16'hfe05;
			16'hfa99: y = 16'hfe05;
			16'hfa9a: y = 16'hfe05;
			16'hfa9b: y = 16'hfe05;
			16'hfa9c: y = 16'hfe05;
			16'hfa9d: y = 16'hfe05;
			16'hfa9e: y = 16'hfe05;
			16'hfa9f: y = 16'hfe05;
			16'hfaa0: y = 16'hfe05;
			16'hfaa1: y = 16'hfe05;
			16'hfaa2: y = 16'hfe05;
			16'hfaa3: y = 16'hfe05;
			16'hfaa4: y = 16'hfe05;
			16'hfaa5: y = 16'hfe05;
			16'hfaa6: y = 16'hfe05;
			16'hfaa7: y = 16'hfe05;
			16'hfaa8: y = 16'hfe05;
			16'hfaa9: y = 16'hfe05;
			16'hfaaa: y = 16'hfe05;
			16'hfaab: y = 16'hfe05;
			16'hfaac: y = 16'hfe05;
			16'hfaad: y = 16'hfe05;
			16'hfaae: y = 16'hfe05;
			16'hfaaf: y = 16'hfe06;
			16'hfab0: y = 16'hfe06;
			16'hfab1: y = 16'hfe06;
			16'hfab2: y = 16'hfe06;
			16'hfab3: y = 16'hfe06;
			16'hfab4: y = 16'hfe06;
			16'hfab5: y = 16'hfe06;
			16'hfab6: y = 16'hfe06;
			16'hfab7: y = 16'hfe06;
			16'hfab8: y = 16'hfe06;
			16'hfab9: y = 16'hfe06;
			16'hfaba: y = 16'hfe06;
			16'hfabb: y = 16'hfe06;
			16'hfabc: y = 16'hfe06;
			16'hfabd: y = 16'hfe06;
			16'hfabe: y = 16'hfe06;
			16'hfabf: y = 16'hfe06;
			16'hfac0: y = 16'hfe06;
			16'hfac1: y = 16'hfe06;
			16'hfac2: y = 16'hfe06;
			16'hfac3: y = 16'hfe06;
			16'hfac4: y = 16'hfe06;
			16'hfac5: y = 16'hfe06;
			16'hfac6: y = 16'hfe06;
			16'hfac7: y = 16'hfe06;
			16'hfac8: y = 16'hfe06;
			16'hfac9: y = 16'hfe06;
			16'hfaca: y = 16'hfe06;
			16'hfacb: y = 16'hfe06;
			16'hfacc: y = 16'hfe06;
			16'hfacd: y = 16'hfe06;
			16'hface: y = 16'hfe06;
			16'hfacf: y = 16'hfe06;
			16'hfad0: y = 16'hfe06;
			16'hfad1: y = 16'hfe06;
			16'hfad2: y = 16'hfe06;
			16'hfad3: y = 16'hfe06;
			16'hfad4: y = 16'hfe06;
			16'hfad5: y = 16'hfe06;
			16'hfad6: y = 16'hfe06;
			16'hfad7: y = 16'hfe06;
			16'hfad8: y = 16'hfe06;
			16'hfad9: y = 16'hfe06;
			16'hfada: y = 16'hfe06;
			16'hfadb: y = 16'hfe06;
			16'hfadc: y = 16'hfe06;
			16'hfadd: y = 16'hfe06;
			16'hfade: y = 16'hfe07;
			16'hfadf: y = 16'hfe07;
			16'hfae0: y = 16'hfe07;
			16'hfae1: y = 16'hfe07;
			16'hfae2: y = 16'hfe07;
			16'hfae3: y = 16'hfe07;
			16'hfae4: y = 16'hfe07;
			16'hfae5: y = 16'hfe07;
			16'hfae6: y = 16'hfe07;
			16'hfae7: y = 16'hfe07;
			16'hfae8: y = 16'hfe07;
			16'hfae9: y = 16'hfe07;
			16'hfaea: y = 16'hfe07;
			16'hfaeb: y = 16'hfe07;
			16'hfaec: y = 16'hfe07;
			16'hfaed: y = 16'hfe07;
			16'hfaee: y = 16'hfe07;
			16'hfaef: y = 16'hfe07;
			16'hfaf0: y = 16'hfe07;
			16'hfaf1: y = 16'hfe07;
			16'hfaf2: y = 16'hfe07;
			16'hfaf3: y = 16'hfe07;
			16'hfaf4: y = 16'hfe07;
			16'hfaf5: y = 16'hfe07;
			16'hfaf6: y = 16'hfe07;
			16'hfaf7: y = 16'hfe07;
			16'hfaf8: y = 16'hfe07;
			16'hfaf9: y = 16'hfe07;
			16'hfafa: y = 16'hfe07;
			16'hfafb: y = 16'hfe07;
			16'hfafc: y = 16'hfe07;
			16'hfafd: y = 16'hfe07;
			16'hfafe: y = 16'hfe07;
			16'hfaff: y = 16'hfe07;
			16'hfb00: y = 16'hfe07;
			16'hfb01: y = 16'hfe07;
			16'hfb02: y = 16'hfe07;
			16'hfb03: y = 16'hfe07;
			16'hfb04: y = 16'hfe07;
			16'hfb05: y = 16'hfe07;
			16'hfb06: y = 16'hfe08;
			16'hfb07: y = 16'hfe08;
			16'hfb08: y = 16'hfe08;
			16'hfb09: y = 16'hfe08;
			16'hfb0a: y = 16'hfe08;
			16'hfb0b: y = 16'hfe08;
			16'hfb0c: y = 16'hfe08;
			16'hfb0d: y = 16'hfe08;
			16'hfb0e: y = 16'hfe08;
			16'hfb0f: y = 16'hfe08;
			16'hfb10: y = 16'hfe08;
			16'hfb11: y = 16'hfe08;
			16'hfb12: y = 16'hfe08;
			16'hfb13: y = 16'hfe08;
			16'hfb14: y = 16'hfe08;
			16'hfb15: y = 16'hfe08;
			16'hfb16: y = 16'hfe08;
			16'hfb17: y = 16'hfe08;
			16'hfb18: y = 16'hfe08;
			16'hfb19: y = 16'hfe08;
			16'hfb1a: y = 16'hfe08;
			16'hfb1b: y = 16'hfe08;
			16'hfb1c: y = 16'hfe08;
			16'hfb1d: y = 16'hfe08;
			16'hfb1e: y = 16'hfe08;
			16'hfb1f: y = 16'hfe08;
			16'hfb20: y = 16'hfe08;
			16'hfb21: y = 16'hfe08;
			16'hfb22: y = 16'hfe08;
			16'hfb23: y = 16'hfe08;
			16'hfb24: y = 16'hfe08;
			16'hfb25: y = 16'hfe08;
			16'hfb26: y = 16'hfe08;
			16'hfb27: y = 16'hfe08;
			16'hfb28: y = 16'hfe09;
			16'hfb29: y = 16'hfe09;
			16'hfb2a: y = 16'hfe09;
			16'hfb2b: y = 16'hfe09;
			16'hfb2c: y = 16'hfe09;
			16'hfb2d: y = 16'hfe09;
			16'hfb2e: y = 16'hfe09;
			16'hfb2f: y = 16'hfe09;
			16'hfb30: y = 16'hfe09;
			16'hfb31: y = 16'hfe09;
			16'hfb32: y = 16'hfe09;
			16'hfb33: y = 16'hfe09;
			16'hfb34: y = 16'hfe09;
			16'hfb35: y = 16'hfe09;
			16'hfb36: y = 16'hfe09;
			16'hfb37: y = 16'hfe09;
			16'hfb38: y = 16'hfe09;
			16'hfb39: y = 16'hfe09;
			16'hfb3a: y = 16'hfe09;
			16'hfb3b: y = 16'hfe09;
			16'hfb3c: y = 16'hfe09;
			16'hfb3d: y = 16'hfe09;
			16'hfb3e: y = 16'hfe09;
			16'hfb3f: y = 16'hfe09;
			16'hfb40: y = 16'hfe09;
			16'hfb41: y = 16'hfe09;
			16'hfb42: y = 16'hfe09;
			16'hfb43: y = 16'hfe09;
			16'hfb44: y = 16'hfe09;
			16'hfb45: y = 16'hfe09;
			16'hfb46: y = 16'hfe09;
			16'hfb47: y = 16'hfe0a;
			16'hfb48: y = 16'hfe0a;
			16'hfb49: y = 16'hfe0a;
			16'hfb4a: y = 16'hfe0a;
			16'hfb4b: y = 16'hfe0a;
			16'hfb4c: y = 16'hfe0a;
			16'hfb4d: y = 16'hfe0a;
			16'hfb4e: y = 16'hfe0a;
			16'hfb4f: y = 16'hfe0a;
			16'hfb50: y = 16'hfe0a;
			16'hfb51: y = 16'hfe0a;
			16'hfb52: y = 16'hfe0a;
			16'hfb53: y = 16'hfe0a;
			16'hfb54: y = 16'hfe0a;
			16'hfb55: y = 16'hfe0a;
			16'hfb56: y = 16'hfe0a;
			16'hfb57: y = 16'hfe0a;
			16'hfb58: y = 16'hfe0a;
			16'hfb59: y = 16'hfe0a;
			16'hfb5a: y = 16'hfe0a;
			16'hfb5b: y = 16'hfe0a;
			16'hfb5c: y = 16'hfe0a;
			16'hfb5d: y = 16'hfe0a;
			16'hfb5e: y = 16'hfe0a;
			16'hfb5f: y = 16'hfe0a;
			16'hfb60: y = 16'hfe0a;
			16'hfb61: y = 16'hfe0a;
			16'hfb62: y = 16'hfe0b;
			16'hfb63: y = 16'hfe0b;
			16'hfb64: y = 16'hfe0b;
			16'hfb65: y = 16'hfe0b;
			16'hfb66: y = 16'hfe0b;
			16'hfb67: y = 16'hfe0b;
			16'hfb68: y = 16'hfe0b;
			16'hfb69: y = 16'hfe0b;
			16'hfb6a: y = 16'hfe0b;
			16'hfb6b: y = 16'hfe0b;
			16'hfb6c: y = 16'hfe0b;
			16'hfb6d: y = 16'hfe0b;
			16'hfb6e: y = 16'hfe0b;
			16'hfb6f: y = 16'hfe0b;
			16'hfb70: y = 16'hfe0b;
			16'hfb71: y = 16'hfe0b;
			16'hfb72: y = 16'hfe0b;
			16'hfb73: y = 16'hfe0b;
			16'hfb74: y = 16'hfe0b;
			16'hfb75: y = 16'hfe0b;
			16'hfb76: y = 16'hfe0b;
			16'hfb77: y = 16'hfe0b;
			16'hfb78: y = 16'hfe0b;
			16'hfb79: y = 16'hfe0b;
			16'hfb7a: y = 16'hfe0b;
			16'hfb7b: y = 16'hfe0c;
			16'hfb7c: y = 16'hfe0c;
			16'hfb7d: y = 16'hfe0c;
			16'hfb7e: y = 16'hfe0c;
			16'hfb7f: y = 16'hfe0c;
			16'hfb80: y = 16'hfe0c;
			16'hfb81: y = 16'hfe0c;
			16'hfb82: y = 16'hfe0c;
			16'hfb83: y = 16'hfe0c;
			16'hfb84: y = 16'hfe0c;
			16'hfb85: y = 16'hfe0c;
			16'hfb86: y = 16'hfe0c;
			16'hfb87: y = 16'hfe0c;
			16'hfb88: y = 16'hfe0c;
			16'hfb89: y = 16'hfe0c;
			16'hfb8a: y = 16'hfe0c;
			16'hfb8b: y = 16'hfe0c;
			16'hfb8c: y = 16'hfe0c;
			16'hfb8d: y = 16'hfe0c;
			16'hfb8e: y = 16'hfe0c;
			16'hfb8f: y = 16'hfe0c;
			16'hfb90: y = 16'hfe0c;
			16'hfb91: y = 16'hfe0d;
			16'hfb92: y = 16'hfe0d;
			16'hfb93: y = 16'hfe0d;
			16'hfb94: y = 16'hfe0d;
			16'hfb95: y = 16'hfe0d;
			16'hfb96: y = 16'hfe0d;
			16'hfb97: y = 16'hfe0d;
			16'hfb98: y = 16'hfe0d;
			16'hfb99: y = 16'hfe0d;
			16'hfb9a: y = 16'hfe0d;
			16'hfb9b: y = 16'hfe0d;
			16'hfb9c: y = 16'hfe0d;
			16'hfb9d: y = 16'hfe0d;
			16'hfb9e: y = 16'hfe0d;
			16'hfb9f: y = 16'hfe0d;
			16'hfba0: y = 16'hfe0d;
			16'hfba1: y = 16'hfe0d;
			16'hfba2: y = 16'hfe0d;
			16'hfba3: y = 16'hfe0d;
			16'hfba4: y = 16'hfe0d;
			16'hfba5: y = 16'hfe0d;
			16'hfba6: y = 16'hfe0e;
			16'hfba7: y = 16'hfe0e;
			16'hfba8: y = 16'hfe0e;
			16'hfba9: y = 16'hfe0e;
			16'hfbaa: y = 16'hfe0e;
			16'hfbab: y = 16'hfe0e;
			16'hfbac: y = 16'hfe0e;
			16'hfbad: y = 16'hfe0e;
			16'hfbae: y = 16'hfe0e;
			16'hfbaf: y = 16'hfe0e;
			16'hfbb0: y = 16'hfe0e;
			16'hfbb1: y = 16'hfe0e;
			16'hfbb2: y = 16'hfe0e;
			16'hfbb3: y = 16'hfe0e;
			16'hfbb4: y = 16'hfe0e;
			16'hfbb5: y = 16'hfe0e;
			16'hfbb6: y = 16'hfe0e;
			16'hfbb7: y = 16'hfe0e;
			16'hfbb8: y = 16'hfe0e;
			16'hfbb9: y = 16'hfe0f;
			16'hfbba: y = 16'hfe0f;
			16'hfbbb: y = 16'hfe0f;
			16'hfbbc: y = 16'hfe0f;
			16'hfbbd: y = 16'hfe0f;
			16'hfbbe: y = 16'hfe0f;
			16'hfbbf: y = 16'hfe0f;
			16'hfbc0: y = 16'hfe0f;
			16'hfbc1: y = 16'hfe0f;
			16'hfbc2: y = 16'hfe0f;
			16'hfbc3: y = 16'hfe0f;
			16'hfbc4: y = 16'hfe0f;
			16'hfbc5: y = 16'hfe0f;
			16'hfbc6: y = 16'hfe0f;
			16'hfbc7: y = 16'hfe0f;
			16'hfbc8: y = 16'hfe0f;
			16'hfbc9: y = 16'hfe0f;
			16'hfbca: y = 16'hfe0f;
			16'hfbcb: y = 16'hfe10;
			16'hfbcc: y = 16'hfe10;
			16'hfbcd: y = 16'hfe10;
			16'hfbce: y = 16'hfe10;
			16'hfbcf: y = 16'hfe10;
			16'hfbd0: y = 16'hfe10;
			16'hfbd1: y = 16'hfe10;
			16'hfbd2: y = 16'hfe10;
			16'hfbd3: y = 16'hfe10;
			16'hfbd4: y = 16'hfe10;
			16'hfbd5: y = 16'hfe10;
			16'hfbd6: y = 16'hfe10;
			16'hfbd7: y = 16'hfe10;
			16'hfbd8: y = 16'hfe10;
			16'hfbd9: y = 16'hfe10;
			16'hfbda: y = 16'hfe10;
			16'hfbdb: y = 16'hfe10;
			16'hfbdc: y = 16'hfe11;
			16'hfbdd: y = 16'hfe11;
			16'hfbde: y = 16'hfe11;
			16'hfbdf: y = 16'hfe11;
			16'hfbe0: y = 16'hfe11;
			16'hfbe1: y = 16'hfe11;
			16'hfbe2: y = 16'hfe11;
			16'hfbe3: y = 16'hfe11;
			16'hfbe4: y = 16'hfe11;
			16'hfbe5: y = 16'hfe11;
			16'hfbe6: y = 16'hfe11;
			16'hfbe7: y = 16'hfe11;
			16'hfbe8: y = 16'hfe11;
			16'hfbe9: y = 16'hfe11;
			16'hfbea: y = 16'hfe11;
			16'hfbeb: y = 16'hfe11;
			16'hfbec: y = 16'hfe12;
			16'hfbed: y = 16'hfe12;
			16'hfbee: y = 16'hfe12;
			16'hfbef: y = 16'hfe12;
			16'hfbf0: y = 16'hfe12;
			16'hfbf1: y = 16'hfe12;
			16'hfbf2: y = 16'hfe12;
			16'hfbf3: y = 16'hfe12;
			16'hfbf4: y = 16'hfe12;
			16'hfbf5: y = 16'hfe12;
			16'hfbf6: y = 16'hfe12;
			16'hfbf7: y = 16'hfe12;
			16'hfbf8: y = 16'hfe12;
			16'hfbf9: y = 16'hfe12;
			16'hfbfa: y = 16'hfe12;
			16'hfbfb: y = 16'hfe13;
			16'hfbfc: y = 16'hfe13;
			16'hfbfd: y = 16'hfe13;
			16'hfbfe: y = 16'hfe13;
			16'hfbff: y = 16'hfe13;
			16'hfc00: y = 16'hfe13;
			16'hfc01: y = 16'hfe13;
			16'hfc02: y = 16'hfe13;
			16'hfc03: y = 16'hfe13;
			16'hfc04: y = 16'hfe13;
			16'hfc05: y = 16'hfe13;
			16'hfc06: y = 16'hfe13;
			16'hfc07: y = 16'hfe13;
			16'hfc08: y = 16'hfe13;
			16'hfc09: y = 16'hfe14;
			16'hfc0a: y = 16'hfe14;
			16'hfc0b: y = 16'hfe14;
			16'hfc0c: y = 16'hfe14;
			16'hfc0d: y = 16'hfe14;
			16'hfc0e: y = 16'hfe14;
			16'hfc0f: y = 16'hfe14;
			16'hfc10: y = 16'hfe14;
			16'hfc11: y = 16'hfe14;
			16'hfc12: y = 16'hfe14;
			16'hfc13: y = 16'hfe14;
			16'hfc14: y = 16'hfe14;
			16'hfc15: y = 16'hfe14;
			16'hfc16: y = 16'hfe15;
			16'hfc17: y = 16'hfe15;
			16'hfc18: y = 16'hfe15;
			16'hfc19: y = 16'hfe15;
			16'hfc1a: y = 16'hfe15;
			16'hfc1b: y = 16'hfe15;
			16'hfc1c: y = 16'hfe15;
			16'hfc1d: y = 16'hfe15;
			16'hfc1e: y = 16'hfe15;
			16'hfc1f: y = 16'hfe15;
			16'hfc20: y = 16'hfe15;
			16'hfc21: y = 16'hfe15;
			16'hfc22: y = 16'hfe15;
			16'hfc23: y = 16'hfe16;
			16'hfc24: y = 16'hfe16;
			16'hfc25: y = 16'hfe16;
			16'hfc26: y = 16'hfe16;
			16'hfc27: y = 16'hfe16;
			16'hfc28: y = 16'hfe16;
			16'hfc29: y = 16'hfe16;
			16'hfc2a: y = 16'hfe16;
			16'hfc2b: y = 16'hfe16;
			16'hfc2c: y = 16'hfe16;
			16'hfc2d: y = 16'hfe16;
			16'hfc2e: y = 16'hfe16;
			16'hfc2f: y = 16'hfe17;
			16'hfc30: y = 16'hfe17;
			16'hfc31: y = 16'hfe17;
			16'hfc32: y = 16'hfe17;
			16'hfc33: y = 16'hfe17;
			16'hfc34: y = 16'hfe17;
			16'hfc35: y = 16'hfe17;
			16'hfc36: y = 16'hfe17;
			16'hfc37: y = 16'hfe17;
			16'hfc38: y = 16'hfe17;
			16'hfc39: y = 16'hfe17;
			16'hfc3a: y = 16'hfe17;
			16'hfc3b: y = 16'hfe18;
			16'hfc3c: y = 16'hfe18;
			16'hfc3d: y = 16'hfe18;
			16'hfc3e: y = 16'hfe18;
			16'hfc3f: y = 16'hfe18;
			16'hfc40: y = 16'hfe18;
			16'hfc41: y = 16'hfe18;
			16'hfc42: y = 16'hfe18;
			16'hfc43: y = 16'hfe18;
			16'hfc44: y = 16'hfe18;
			16'hfc45: y = 16'hfe18;
			16'hfc46: y = 16'hfe19;
			16'hfc47: y = 16'hfe19;
			16'hfc48: y = 16'hfe19;
			16'hfc49: y = 16'hfe19;
			16'hfc4a: y = 16'hfe19;
			16'hfc4b: y = 16'hfe19;
			16'hfc4c: y = 16'hfe19;
			16'hfc4d: y = 16'hfe19;
			16'hfc4e: y = 16'hfe19;
			16'hfc4f: y = 16'hfe19;
			16'hfc50: y = 16'hfe1a;
			16'hfc51: y = 16'hfe1a;
			16'hfc52: y = 16'hfe1a;
			16'hfc53: y = 16'hfe1a;
			16'hfc54: y = 16'hfe1a;
			16'hfc55: y = 16'hfe1a;
			16'hfc56: y = 16'hfe1a;
			16'hfc57: y = 16'hfe1a;
			16'hfc58: y = 16'hfe1a;
			16'hfc59: y = 16'hfe1a;
			16'hfc5a: y = 16'hfe1a;
			16'hfc5b: y = 16'hfe1b;
			16'hfc5c: y = 16'hfe1b;
			16'hfc5d: y = 16'hfe1b;
			16'hfc5e: y = 16'hfe1b;
			16'hfc5f: y = 16'hfe1b;
			16'hfc60: y = 16'hfe1b;
			16'hfc61: y = 16'hfe1b;
			16'hfc62: y = 16'hfe1b;
			16'hfc63: y = 16'hfe1b;
			16'hfc64: y = 16'hfe1b;
			16'hfc65: y = 16'hfe1c;
			16'hfc66: y = 16'hfe1c;
			16'hfc67: y = 16'hfe1c;
			16'hfc68: y = 16'hfe1c;
			16'hfc69: y = 16'hfe1c;
			16'hfc6a: y = 16'hfe1c;
			16'hfc6b: y = 16'hfe1c;
			16'hfc6c: y = 16'hfe1c;
			16'hfc6d: y = 16'hfe1c;
			16'hfc6e: y = 16'hfe1d;
			16'hfc6f: y = 16'hfe1d;
			16'hfc70: y = 16'hfe1d;
			16'hfc71: y = 16'hfe1d;
			16'hfc72: y = 16'hfe1d;
			16'hfc73: y = 16'hfe1d;
			16'hfc74: y = 16'hfe1d;
			16'hfc75: y = 16'hfe1d;
			16'hfc76: y = 16'hfe1d;
			16'hfc77: y = 16'hfe1e;
			16'hfc78: y = 16'hfe1e;
			16'hfc79: y = 16'hfe1e;
			16'hfc7a: y = 16'hfe1e;
			16'hfc7b: y = 16'hfe1e;
			16'hfc7c: y = 16'hfe1e;
			16'hfc7d: y = 16'hfe1e;
			16'hfc7e: y = 16'hfe1e;
			16'hfc7f: y = 16'hfe1e;
			16'hfc80: y = 16'hfe1f;
			16'hfc81: y = 16'hfe1f;
			16'hfc82: y = 16'hfe1f;
			16'hfc83: y = 16'hfe1f;
			16'hfc84: y = 16'hfe1f;
			16'hfc85: y = 16'hfe1f;
			16'hfc86: y = 16'hfe1f;
			16'hfc87: y = 16'hfe1f;
			16'hfc88: y = 16'hfe1f;
			16'hfc89: y = 16'hfe20;
			16'hfc8a: y = 16'hfe20;
			16'hfc8b: y = 16'hfe20;
			16'hfc8c: y = 16'hfe20;
			16'hfc8d: y = 16'hfe20;
			16'hfc8e: y = 16'hfe20;
			16'hfc8f: y = 16'hfe20;
			16'hfc90: y = 16'hfe20;
			16'hfc91: y = 16'hfe21;
			16'hfc92: y = 16'hfe21;
			16'hfc93: y = 16'hfe21;
			16'hfc94: y = 16'hfe21;
			16'hfc95: y = 16'hfe21;
			16'hfc96: y = 16'hfe21;
			16'hfc97: y = 16'hfe21;
			16'hfc98: y = 16'hfe21;
			16'hfc99: y = 16'hfe21;
			16'hfc9a: y = 16'hfe22;
			16'hfc9b: y = 16'hfe22;
			16'hfc9c: y = 16'hfe22;
			16'hfc9d: y = 16'hfe22;
			16'hfc9e: y = 16'hfe22;
			16'hfc9f: y = 16'hfe22;
			16'hfca0: y = 16'hfe22;
			16'hfca1: y = 16'hfe23;
			16'hfca2: y = 16'hfe23;
			16'hfca3: y = 16'hfe23;
			16'hfca4: y = 16'hfe23;
			16'hfca5: y = 16'hfe23;
			16'hfca6: y = 16'hfe23;
			16'hfca7: y = 16'hfe23;
			16'hfca8: y = 16'hfe23;
			16'hfca9: y = 16'hfe24;
			16'hfcaa: y = 16'hfe24;
			16'hfcab: y = 16'hfe24;
			16'hfcac: y = 16'hfe24;
			16'hfcad: y = 16'hfe24;
			16'hfcae: y = 16'hfe24;
			16'hfcaf: y = 16'hfe24;
			16'hfcb0: y = 16'hfe24;
			16'hfcb1: y = 16'hfe25;
			16'hfcb2: y = 16'hfe25;
			16'hfcb3: y = 16'hfe25;
			16'hfcb4: y = 16'hfe25;
			16'hfcb5: y = 16'hfe25;
			16'hfcb6: y = 16'hfe25;
			16'hfcb7: y = 16'hfe25;
			16'hfcb8: y = 16'hfe26;
			16'hfcb9: y = 16'hfe26;
			16'hfcba: y = 16'hfe26;
			16'hfcbb: y = 16'hfe26;
			16'hfcbc: y = 16'hfe26;
			16'hfcbd: y = 16'hfe26;
			16'hfcbe: y = 16'hfe26;
			16'hfcbf: y = 16'hfe27;
			16'hfcc0: y = 16'hfe27;
			16'hfcc1: y = 16'hfe27;
			16'hfcc2: y = 16'hfe27;
			16'hfcc3: y = 16'hfe27;
			16'hfcc4: y = 16'hfe27;
			16'hfcc5: y = 16'hfe27;
			16'hfcc6: y = 16'hfe28;
			16'hfcc7: y = 16'hfe28;
			16'hfcc8: y = 16'hfe28;
			16'hfcc9: y = 16'hfe28;
			16'hfcca: y = 16'hfe28;
			16'hfccb: y = 16'hfe28;
			16'hfccc: y = 16'hfe28;
			16'hfccd: y = 16'hfe29;
			16'hfcce: y = 16'hfe29;
			16'hfccf: y = 16'hfe29;
			16'hfcd0: y = 16'hfe29;
			16'hfcd1: y = 16'hfe29;
			16'hfcd2: y = 16'hfe29;
			16'hfcd3: y = 16'hfe2a;
			16'hfcd4: y = 16'hfe2a;
			16'hfcd5: y = 16'hfe2a;
			16'hfcd6: y = 16'hfe2a;
			16'hfcd7: y = 16'hfe2a;
			16'hfcd8: y = 16'hfe2a;
			16'hfcd9: y = 16'hfe2a;
			16'hfcda: y = 16'hfe2b;
			16'hfcdb: y = 16'hfe2b;
			16'hfcdc: y = 16'hfe2b;
			16'hfcdd: y = 16'hfe2b;
			16'hfcde: y = 16'hfe2b;
			16'hfcdf: y = 16'hfe2b;
			16'hfce0: y = 16'hfe2c;
			16'hfce1: y = 16'hfe2c;
			16'hfce2: y = 16'hfe2c;
			16'hfce3: y = 16'hfe2c;
			16'hfce4: y = 16'hfe2c;
			16'hfce5: y = 16'hfe2c;
			16'hfce6: y = 16'hfe2d;
			16'hfce7: y = 16'hfe2d;
			16'hfce8: y = 16'hfe2d;
			16'hfce9: y = 16'hfe2d;
			16'hfcea: y = 16'hfe2d;
			16'hfceb: y = 16'hfe2d;
			16'hfcec: y = 16'hfe2e;
			16'hfced: y = 16'hfe2e;
			16'hfcee: y = 16'hfe2e;
			16'hfcef: y = 16'hfe2e;
			16'hfcf0: y = 16'hfe2e;
			16'hfcf1: y = 16'hfe2e;
			16'hfcf2: y = 16'hfe2f;
			16'hfcf3: y = 16'hfe2f;
			16'hfcf4: y = 16'hfe2f;
			16'hfcf5: y = 16'hfe2f;
			16'hfcf6: y = 16'hfe2f;
			16'hfcf7: y = 16'hfe2f;
			16'hfcf8: y = 16'hfe30;
			16'hfcf9: y = 16'hfe30;
			16'hfcfa: y = 16'hfe30;
			16'hfcfb: y = 16'hfe30;
			16'hfcfc: y = 16'hfe30;
			16'hfcfd: y = 16'hfe31;
			16'hfcfe: y = 16'hfe31;
			16'hfcff: y = 16'hfe31;
			16'hfd00: y = 16'hfe31;
			16'hfd01: y = 16'hfe31;
			16'hfd02: y = 16'hfe31;
			16'hfd03: y = 16'hfe32;
			16'hfd04: y = 16'hfe32;
			16'hfd05: y = 16'hfe32;
			16'hfd06: y = 16'hfe32;
			16'hfd07: y = 16'hfe32;
			16'hfd08: y = 16'hfe33;
			16'hfd09: y = 16'hfe33;
			16'hfd0a: y = 16'hfe33;
			16'hfd0b: y = 16'hfe33;
			16'hfd0c: y = 16'hfe33;
			16'hfd0d: y = 16'hfe33;
			16'hfd0e: y = 16'hfe34;
			16'hfd0f: y = 16'hfe34;
			16'hfd10: y = 16'hfe34;
			16'hfd11: y = 16'hfe34;
			16'hfd12: y = 16'hfe34;
			16'hfd13: y = 16'hfe35;
			16'hfd14: y = 16'hfe35;
			16'hfd15: y = 16'hfe35;
			16'hfd16: y = 16'hfe35;
			16'hfd17: y = 16'hfe35;
			16'hfd18: y = 16'hfe36;
			16'hfd19: y = 16'hfe36;
			16'hfd1a: y = 16'hfe36;
			16'hfd1b: y = 16'hfe36;
			16'hfd1c: y = 16'hfe36;
			16'hfd1d: y = 16'hfe37;
			16'hfd1e: y = 16'hfe37;
			16'hfd1f: y = 16'hfe37;
			16'hfd20: y = 16'hfe37;
			16'hfd21: y = 16'hfe37;
			16'hfd22: y = 16'hfe38;
			16'hfd23: y = 16'hfe38;
			16'hfd24: y = 16'hfe38;
			16'hfd25: y = 16'hfe38;
			16'hfd26: y = 16'hfe38;
			16'hfd27: y = 16'hfe39;
			16'hfd28: y = 16'hfe39;
			16'hfd29: y = 16'hfe39;
			16'hfd2a: y = 16'hfe39;
			16'hfd2b: y = 16'hfe39;
			16'hfd2c: y = 16'hfe3a;
			16'hfd2d: y = 16'hfe3a;
			16'hfd2e: y = 16'hfe3a;
			16'hfd2f: y = 16'hfe3a;
			16'hfd30: y = 16'hfe3b;
			16'hfd31: y = 16'hfe3b;
			16'hfd32: y = 16'hfe3b;
			16'hfd33: y = 16'hfe3b;
			16'hfd34: y = 16'hfe3b;
			16'hfd35: y = 16'hfe3c;
			16'hfd36: y = 16'hfe3c;
			16'hfd37: y = 16'hfe3c;
			16'hfd38: y = 16'hfe3c;
			16'hfd39: y = 16'hfe3c;
			16'hfd3a: y = 16'hfe3d;
			16'hfd3b: y = 16'hfe3d;
			16'hfd3c: y = 16'hfe3d;
			16'hfd3d: y = 16'hfe3d;
			16'hfd3e: y = 16'hfe3e;
			16'hfd3f: y = 16'hfe3e;
			16'hfd40: y = 16'hfe3e;
			16'hfd41: y = 16'hfe3e;
			16'hfd42: y = 16'hfe3e;
			16'hfd43: y = 16'hfe3f;
			16'hfd44: y = 16'hfe3f;
			16'hfd45: y = 16'hfe3f;
			16'hfd46: y = 16'hfe3f;
			16'hfd47: y = 16'hfe40;
			16'hfd48: y = 16'hfe40;
			16'hfd49: y = 16'hfe40;
			16'hfd4a: y = 16'hfe40;
			16'hfd4b: y = 16'hfe41;
			16'hfd4c: y = 16'hfe41;
			16'hfd4d: y = 16'hfe41;
			16'hfd4e: y = 16'hfe41;
			16'hfd4f: y = 16'hfe42;
			16'hfd50: y = 16'hfe42;
			16'hfd51: y = 16'hfe42;
			16'hfd52: y = 16'hfe42;
			16'hfd53: y = 16'hfe42;
			16'hfd54: y = 16'hfe43;
			16'hfd55: y = 16'hfe43;
			16'hfd56: y = 16'hfe43;
			16'hfd57: y = 16'hfe43;
			16'hfd58: y = 16'hfe44;
			16'hfd59: y = 16'hfe44;
			16'hfd5a: y = 16'hfe44;
			16'hfd5b: y = 16'hfe44;
			16'hfd5c: y = 16'hfe45;
			16'hfd5d: y = 16'hfe45;
			16'hfd5e: y = 16'hfe45;
			16'hfd5f: y = 16'hfe45;
			16'hfd60: y = 16'hfe46;
			16'hfd61: y = 16'hfe46;
			16'hfd62: y = 16'hfe46;
			16'hfd63: y = 16'hfe46;
			16'hfd64: y = 16'hfe47;
			16'hfd65: y = 16'hfe47;
			16'hfd66: y = 16'hfe47;
			16'hfd67: y = 16'hfe47;
			16'hfd68: y = 16'hfe48;
			16'hfd69: y = 16'hfe48;
			16'hfd6a: y = 16'hfe48;
			16'hfd6b: y = 16'hfe48;
			16'hfd6c: y = 16'hfe49;
			16'hfd6d: y = 16'hfe49;
			16'hfd6e: y = 16'hfe49;
			16'hfd6f: y = 16'hfe4a;
			16'hfd70: y = 16'hfe4a;
			16'hfd71: y = 16'hfe4a;
			16'hfd72: y = 16'hfe4a;
			16'hfd73: y = 16'hfe4b;
			16'hfd74: y = 16'hfe4b;
			16'hfd75: y = 16'hfe4b;
			16'hfd76: y = 16'hfe4b;
			16'hfd77: y = 16'hfe4c;
			16'hfd78: y = 16'hfe4c;
			16'hfd79: y = 16'hfe4c;
			16'hfd7a: y = 16'hfe4d;
			16'hfd7b: y = 16'hfe4d;
			16'hfd7c: y = 16'hfe4d;
			16'hfd7d: y = 16'hfe4d;
			16'hfd7e: y = 16'hfe4e;
			16'hfd7f: y = 16'hfe4e;
			16'hfd80: y = 16'hfe4e;
			16'hfd81: y = 16'hfe4e;
			16'hfd82: y = 16'hfe4f;
			16'hfd83: y = 16'hfe4f;
			16'hfd84: y = 16'hfe4f;
			16'hfd85: y = 16'hfe50;
			16'hfd86: y = 16'hfe50;
			16'hfd87: y = 16'hfe50;
			16'hfd88: y = 16'hfe50;
			16'hfd89: y = 16'hfe51;
			16'hfd8a: y = 16'hfe51;
			16'hfd8b: y = 16'hfe51;
			16'hfd8c: y = 16'hfe52;
			16'hfd8d: y = 16'hfe52;
			16'hfd8e: y = 16'hfe52;
			16'hfd8f: y = 16'hfe52;
			16'hfd90: y = 16'hfe53;
			16'hfd91: y = 16'hfe53;
			16'hfd92: y = 16'hfe53;
			16'hfd93: y = 16'hfe54;
			16'hfd94: y = 16'hfe54;
			16'hfd95: y = 16'hfe54;
			16'hfd96: y = 16'hfe55;
			16'hfd97: y = 16'hfe55;
			16'hfd98: y = 16'hfe55;
			16'hfd99: y = 16'hfe55;
			16'hfd9a: y = 16'hfe56;
			16'hfd9b: y = 16'hfe56;
			16'hfd9c: y = 16'hfe56;
			16'hfd9d: y = 16'hfe57;
			16'hfd9e: y = 16'hfe57;
			16'hfd9f: y = 16'hfe57;
			16'hfda0: y = 16'hfe58;
			16'hfda1: y = 16'hfe58;
			16'hfda2: y = 16'hfe58;
			16'hfda3: y = 16'hfe59;
			16'hfda4: y = 16'hfe59;
			16'hfda5: y = 16'hfe59;
			16'hfda6: y = 16'hfe5a;
			16'hfda7: y = 16'hfe5a;
			16'hfda8: y = 16'hfe5a;
			16'hfda9: y = 16'hfe5a;
			16'hfdaa: y = 16'hfe5b;
			16'hfdab: y = 16'hfe5b;
			16'hfdac: y = 16'hfe5b;
			16'hfdad: y = 16'hfe5c;
			16'hfdae: y = 16'hfe5c;
			16'hfdaf: y = 16'hfe5c;
			16'hfdb0: y = 16'hfe5d;
			16'hfdb1: y = 16'hfe5d;
			16'hfdb2: y = 16'hfe5d;
			16'hfdb3: y = 16'hfe5e;
			16'hfdb4: y = 16'hfe5e;
			16'hfdb5: y = 16'hfe5e;
			16'hfdb6: y = 16'hfe5f;
			16'hfdb7: y = 16'hfe5f;
			16'hfdb8: y = 16'hfe5f;
			16'hfdb9: y = 16'hfe60;
			16'hfdba: y = 16'hfe60;
			16'hfdbb: y = 16'hfe60;
			16'hfdbc: y = 16'hfe61;
			16'hfdbd: y = 16'hfe61;
			16'hfdbe: y = 16'hfe61;
			16'hfdbf: y = 16'hfe62;
			16'hfdc0: y = 16'hfe62;
			16'hfdc1: y = 16'hfe62;
			16'hfdc2: y = 16'hfe63;
			16'hfdc3: y = 16'hfe63;
			16'hfdc4: y = 16'hfe64;
			16'hfdc5: y = 16'hfe64;
			16'hfdc6: y = 16'hfe64;
			16'hfdc7: y = 16'hfe65;
			16'hfdc8: y = 16'hfe65;
			16'hfdc9: y = 16'hfe65;
			16'hfdca: y = 16'hfe66;
			16'hfdcb: y = 16'hfe66;
			16'hfdcc: y = 16'hfe66;
			16'hfdcd: y = 16'hfe67;
			16'hfdce: y = 16'hfe67;
			16'hfdcf: y = 16'hfe67;
			16'hfdd0: y = 16'hfe68;
			16'hfdd1: y = 16'hfe68;
			16'hfdd2: y = 16'hfe69;
			16'hfdd3: y = 16'hfe69;
			16'hfdd4: y = 16'hfe69;
			16'hfdd5: y = 16'hfe6a;
			16'hfdd6: y = 16'hfe6a;
			16'hfdd7: y = 16'hfe6a;
			16'hfdd8: y = 16'hfe6b;
			16'hfdd9: y = 16'hfe6b;
			16'hfdda: y = 16'hfe6b;
			16'hfddb: y = 16'hfe6c;
			16'hfddc: y = 16'hfe6c;
			16'hfddd: y = 16'hfe6d;
			16'hfdde: y = 16'hfe6d;
			16'hfddf: y = 16'hfe6d;
			16'hfde0: y = 16'hfe6e;
			16'hfde1: y = 16'hfe6e;
			16'hfde2: y = 16'hfe6f;
			16'hfde3: y = 16'hfe6f;
			16'hfde4: y = 16'hfe6f;
			16'hfde5: y = 16'hfe70;
			16'hfde6: y = 16'hfe70;
			16'hfde7: y = 16'hfe70;
			16'hfde8: y = 16'hfe71;
			16'hfde9: y = 16'hfe71;
			16'hfdea: y = 16'hfe72;
			16'hfdeb: y = 16'hfe72;
			16'hfdec: y = 16'hfe72;
			16'hfded: y = 16'hfe73;
			16'hfdee: y = 16'hfe73;
			16'hfdef: y = 16'hfe74;
			16'hfdf0: y = 16'hfe74;
			16'hfdf1: y = 16'hfe74;
			16'hfdf2: y = 16'hfe75;
			16'hfdf3: y = 16'hfe75;
			16'hfdf4: y = 16'hfe76;
			16'hfdf5: y = 16'hfe76;
			16'hfdf6: y = 16'hfe76;
			16'hfdf7: y = 16'hfe77;
			16'hfdf8: y = 16'hfe77;
			16'hfdf9: y = 16'hfe78;
			16'hfdfa: y = 16'hfe78;
			16'hfdfb: y = 16'hfe78;
			16'hfdfc: y = 16'hfe79;
			16'hfdfd: y = 16'hfe79;
			16'hfdfe: y = 16'hfe7a;
			16'hfdff: y = 16'hfe7a;
			16'hfe00: y = 16'hfe7b;
			16'hfe01: y = 16'hfe7b;
			16'hfe02: y = 16'hfe7b;
			16'hfe03: y = 16'hfe7c;
			16'hfe04: y = 16'hfe7c;
			16'hfe05: y = 16'hfe7d;
			16'hfe06: y = 16'hfe7d;
			16'hfe07: y = 16'hfe7e;
			16'hfe08: y = 16'hfe7e;
			16'hfe09: y = 16'hfe7e;
			16'hfe0a: y = 16'hfe7f;
			16'hfe0b: y = 16'hfe7f;
			16'hfe0c: y = 16'hfe80;
			16'hfe0d: y = 16'hfe80;
			16'hfe0e: y = 16'hfe81;
			16'hfe0f: y = 16'hfe81;
			16'hfe10: y = 16'hfe81;
			16'hfe11: y = 16'hfe82;
			16'hfe12: y = 16'hfe82;
			16'hfe13: y = 16'hfe83;
			16'hfe14: y = 16'hfe83;
			16'hfe15: y = 16'hfe84;
			16'hfe16: y = 16'hfe84;
			16'hfe17: y = 16'hfe85;
			16'hfe18: y = 16'hfe85;
			16'hfe19: y = 16'hfe85;
			16'hfe1a: y = 16'hfe86;
			16'hfe1b: y = 16'hfe86;
			16'hfe1c: y = 16'hfe87;
			16'hfe1d: y = 16'hfe87;
			16'hfe1e: y = 16'hfe88;
			16'hfe1f: y = 16'hfe88;
			16'hfe20: y = 16'hfe89;
			16'hfe21: y = 16'hfe89;
			16'hfe22: y = 16'hfe8a;
			16'hfe23: y = 16'hfe8a;
			16'hfe24: y = 16'hfe8b;
			16'hfe25: y = 16'hfe8b;
			16'hfe26: y = 16'hfe8b;
			16'hfe27: y = 16'hfe8c;
			16'hfe28: y = 16'hfe8c;
			16'hfe29: y = 16'hfe8d;
			16'hfe2a: y = 16'hfe8d;
			16'hfe2b: y = 16'hfe8e;
			16'hfe2c: y = 16'hfe8e;
			16'hfe2d: y = 16'hfe8f;
			16'hfe2e: y = 16'hfe8f;
			16'hfe2f: y = 16'hfe90;
			16'hfe30: y = 16'hfe90;
			16'hfe31: y = 16'hfe91;
			16'hfe32: y = 16'hfe91;
			16'hfe33: y = 16'hfe92;
			16'hfe34: y = 16'hfe92;
			16'hfe35: y = 16'hfe93;
			16'hfe36: y = 16'hfe93;
			16'hfe37: y = 16'hfe94;
			16'hfe38: y = 16'hfe94;
			16'hfe39: y = 16'hfe95;
			16'hfe3a: y = 16'hfe95;
			16'hfe3b: y = 16'hfe96;
			16'hfe3c: y = 16'hfe96;
			16'hfe3d: y = 16'hfe97;
			16'hfe3e: y = 16'hfe97;
			16'hfe3f: y = 16'hfe98;
			16'hfe40: y = 16'hfe98;
			16'hfe41: y = 16'hfe99;
			16'hfe42: y = 16'hfe99;
			16'hfe43: y = 16'hfe9a;
			16'hfe44: y = 16'hfe9a;
			16'hfe45: y = 16'hfe9b;
			16'hfe46: y = 16'hfe9b;
			16'hfe47: y = 16'hfe9c;
			16'hfe48: y = 16'hfe9c;
			16'hfe49: y = 16'hfe9d;
			16'hfe4a: y = 16'hfe9d;
			16'hfe4b: y = 16'hfe9e;
			16'hfe4c: y = 16'hfe9e;
			16'hfe4d: y = 16'hfe9f;
			16'hfe4e: y = 16'hfe9f;
			16'hfe4f: y = 16'hfea0;
			16'hfe50: y = 16'hfea0;
			16'hfe51: y = 16'hfea1;
			16'hfe52: y = 16'hfea1;
			16'hfe53: y = 16'hfea2;
			16'hfe54: y = 16'hfea2;
			16'hfe55: y = 16'hfea3;
			16'hfe56: y = 16'hfea4;
			16'hfe57: y = 16'hfea4;
			16'hfe58: y = 16'hfea5;
			16'hfe59: y = 16'hfea5;
			16'hfe5a: y = 16'hfea6;
			16'hfe5b: y = 16'hfea6;
			16'hfe5c: y = 16'hfea7;
			16'hfe5d: y = 16'hfea7;
			16'hfe5e: y = 16'hfea8;
			16'hfe5f: y = 16'hfea8;
			16'hfe60: y = 16'hfea9;
			16'hfe61: y = 16'hfeaa;
			16'hfe62: y = 16'hfeaa;
			16'hfe63: y = 16'hfeab;
			16'hfe64: y = 16'hfeab;
			16'hfe65: y = 16'hfeac;
			16'hfe66: y = 16'hfeac;
			16'hfe67: y = 16'hfead;
			16'hfe68: y = 16'hfead;
			16'hfe69: y = 16'hfeae;
			16'hfe6a: y = 16'hfeaf;
			16'hfe6b: y = 16'hfeaf;
			16'hfe6c: y = 16'hfeb0;
			16'hfe6d: y = 16'hfeb0;
			16'hfe6e: y = 16'hfeb1;
			16'hfe6f: y = 16'hfeb1;
			16'hfe70: y = 16'hfeb2;
			16'hfe71: y = 16'hfeb3;
			16'hfe72: y = 16'hfeb3;
			16'hfe73: y = 16'hfeb4;
			16'hfe74: y = 16'hfeb4;
			16'hfe75: y = 16'hfeb5;
			16'hfe76: y = 16'hfeb5;
			16'hfe77: y = 16'hfeb6;
			16'hfe78: y = 16'hfeb7;
			16'hfe79: y = 16'hfeb7;
			16'hfe7a: y = 16'hfeb8;
			16'hfe7b: y = 16'hfeb8;
			16'hfe7c: y = 16'hfeb9;
			16'hfe7d: y = 16'hfeba;
			16'hfe7e: y = 16'hfeba;
			16'hfe7f: y = 16'hfebb;
			16'hfe80: y = 16'hfebb;
			16'hfe81: y = 16'hfebc;
			16'hfe82: y = 16'hfebc;
			16'hfe83: y = 16'hfebd;
			16'hfe84: y = 16'hfebe;
			16'hfe85: y = 16'hfebe;
			16'hfe86: y = 16'hfebf;
			16'hfe87: y = 16'hfec0;
			16'hfe88: y = 16'hfec0;
			16'hfe89: y = 16'hfec1;
			16'hfe8a: y = 16'hfec1;
			16'hfe8b: y = 16'hfec2;
			16'hfe8c: y = 16'hfec3;
			16'hfe8d: y = 16'hfec3;
			16'hfe8e: y = 16'hfec4;
			16'hfe8f: y = 16'hfec4;
			16'hfe90: y = 16'hfec5;
			16'hfe91: y = 16'hfec6;
			16'hfe92: y = 16'hfec6;
			16'hfe93: y = 16'hfec7;
			16'hfe94: y = 16'hfec8;
			16'hfe95: y = 16'hfec8;
			16'hfe96: y = 16'hfec9;
			16'hfe97: y = 16'hfec9;
			16'hfe98: y = 16'hfeca;
			16'hfe99: y = 16'hfecb;
			16'hfe9a: y = 16'hfecb;
			16'hfe9b: y = 16'hfecc;
			16'hfe9c: y = 16'hfecd;
			16'hfe9d: y = 16'hfecd;
			16'hfe9e: y = 16'hfece;
			16'hfe9f: y = 16'hfecf;
			16'hfea0: y = 16'hfecf;
			16'hfea1: y = 16'hfed0;
			16'hfea2: y = 16'hfed0;
			16'hfea3: y = 16'hfed1;
			16'hfea4: y = 16'hfed2;
			16'hfea5: y = 16'hfed2;
			16'hfea6: y = 16'hfed3;
			16'hfea7: y = 16'hfed4;
			16'hfea8: y = 16'hfed4;
			16'hfea9: y = 16'hfed5;
			16'hfeaa: y = 16'hfed6;
			16'hfeab: y = 16'hfed6;
			16'hfeac: y = 16'hfed7;
			16'hfead: y = 16'hfed8;
			16'hfeae: y = 16'hfed8;
			16'hfeaf: y = 16'hfed9;
			16'hfeb0: y = 16'hfeda;
			16'hfeb1: y = 16'hfeda;
			16'hfeb2: y = 16'hfedb;
			16'hfeb3: y = 16'hfedc;
			16'hfeb4: y = 16'hfedc;
			16'hfeb5: y = 16'hfedd;
			16'hfeb6: y = 16'hfede;
			16'hfeb7: y = 16'hfede;
			16'hfeb8: y = 16'hfedf;
			16'hfeb9: y = 16'hfee0;
			16'hfeba: y = 16'hfee0;
			16'hfebb: y = 16'hfee1;
			16'hfebc: y = 16'hfee2;
			16'hfebd: y = 16'hfee2;
			16'hfebe: y = 16'hfee3;
			16'hfebf: y = 16'hfee4;
			16'hfec0: y = 16'hfee5;
			16'hfec1: y = 16'hfee5;
			16'hfec2: y = 16'hfee6;
			16'hfec3: y = 16'hfee7;
			16'hfec4: y = 16'hfee7;
			16'hfec5: y = 16'hfee8;
			16'hfec6: y = 16'hfee9;
			16'hfec7: y = 16'hfee9;
			16'hfec8: y = 16'hfeea;
			16'hfec9: y = 16'hfeeb;
			16'hfeca: y = 16'hfeec;
			16'hfecb: y = 16'hfeec;
			16'hfecc: y = 16'hfeed;
			16'hfecd: y = 16'hfeee;
			16'hfece: y = 16'hfeee;
			16'hfecf: y = 16'hfeef;
			16'hfed0: y = 16'hfef0;
			16'hfed1: y = 16'hfef1;
			16'hfed2: y = 16'hfef1;
			16'hfed3: y = 16'hfef2;
			16'hfed4: y = 16'hfef3;
			16'hfed5: y = 16'hfef3;
			16'hfed6: y = 16'hfef4;
			16'hfed7: y = 16'hfef5;
			16'hfed8: y = 16'hfef6;
			16'hfed9: y = 16'hfef6;
			16'hfeda: y = 16'hfef7;
			16'hfedb: y = 16'hfef8;
			16'hfedc: y = 16'hfef9;
			16'hfedd: y = 16'hfef9;
			16'hfede: y = 16'hfefa;
			16'hfedf: y = 16'hfefb;
			16'hfee0: y = 16'hfefb;
			16'hfee1: y = 16'hfefc;
			16'hfee2: y = 16'hfefd;
			16'hfee3: y = 16'hfefe;
			16'hfee4: y = 16'hfefe;
			16'hfee5: y = 16'hfeff;
			16'hfee6: y = 16'hff00;
			16'hfee7: y = 16'hff01;
			16'hfee8: y = 16'hff01;
			16'hfee9: y = 16'hff02;
			16'hfeea: y = 16'hff03;
			16'hfeeb: y = 16'hff04;
			16'hfeec: y = 16'hff04;
			16'hfeed: y = 16'hff05;
			16'hfeee: y = 16'hff06;
			16'hfeef: y = 16'hff07;
			16'hfef0: y = 16'hff07;
			16'hfef1: y = 16'hff08;
			16'hfef2: y = 16'hff09;
			16'hfef3: y = 16'hff0a;
			16'hfef4: y = 16'hff0b;
			16'hfef5: y = 16'hff0b;
			16'hfef6: y = 16'hff0c;
			16'hfef7: y = 16'hff0d;
			16'hfef8: y = 16'hff0e;
			16'hfef9: y = 16'hff0e;
			16'hfefa: y = 16'hff0f;
			16'hfefb: y = 16'hff10;
			16'hfefc: y = 16'hff11;
			16'hfefd: y = 16'hff12;
			16'hfefe: y = 16'hff12;
			16'hfeff: y = 16'hff13;
			16'hff00: y = 16'hff14;
			16'hff01: y = 16'hff15;
			16'hff02: y = 16'hff15;
			16'hff03: y = 16'hff16;
			16'hff04: y = 16'hff17;
			16'hff05: y = 16'hff18;
			16'hff06: y = 16'hff19;
			16'hff07: y = 16'hff19;
			16'hff08: y = 16'hff1a;
			16'hff09: y = 16'hff1b;
			16'hff0a: y = 16'hff1c;
			16'hff0b: y = 16'hff1d;
			16'hff0c: y = 16'hff1d;
			16'hff0d: y = 16'hff1e;
			16'hff0e: y = 16'hff1f;
			16'hff0f: y = 16'hff20;
			16'hff10: y = 16'hff21;
			16'hff11: y = 16'hff21;
			16'hff12: y = 16'hff22;
			16'hff13: y = 16'hff23;
			16'hff14: y = 16'hff24;
			16'hff15: y = 16'hff25;
			16'hff16: y = 16'hff26;
			16'hff17: y = 16'hff26;
			16'hff18: y = 16'hff27;
			16'hff19: y = 16'hff28;
			16'hff1a: y = 16'hff29;
			16'hff1b: y = 16'hff2a;
			16'hff1c: y = 16'hff2a;
			16'hff1d: y = 16'hff2b;
			16'hff1e: y = 16'hff2c;
			16'hff1f: y = 16'hff2d;
			16'hff20: y = 16'hff2e;
			16'hff21: y = 16'hff2f;
			16'hff22: y = 16'hff2f;
			16'hff23: y = 16'hff30;
			16'hff24: y = 16'hff31;
			16'hff25: y = 16'hff32;
			16'hff26: y = 16'hff33;
			16'hff27: y = 16'hff34;
			16'hff28: y = 16'hff34;
			16'hff29: y = 16'hff35;
			16'hff2a: y = 16'hff36;
			16'hff2b: y = 16'hff37;
			16'hff2c: y = 16'hff38;
			16'hff2d: y = 16'hff39;
			16'hff2e: y = 16'hff3a;
			16'hff2f: y = 16'hff3a;
			16'hff30: y = 16'hff3b;
			16'hff31: y = 16'hff3c;
			16'hff32: y = 16'hff3d;
			16'hff33: y = 16'hff3e;
			16'hff34: y = 16'hff3f;
			16'hff35: y = 16'hff40;
			16'hff36: y = 16'hff40;
			16'hff37: y = 16'hff41;
			16'hff38: y = 16'hff42;
			16'hff39: y = 16'hff43;
			16'hff3a: y = 16'hff44;
			16'hff3b: y = 16'hff45;
			16'hff3c: y = 16'hff46;
			16'hff3d: y = 16'hff46;
			16'hff3e: y = 16'hff47;
			16'hff3f: y = 16'hff48;
			16'hff40: y = 16'hff49;
			16'hff41: y = 16'hff4a;
			16'hff42: y = 16'hff4b;
			16'hff43: y = 16'hff4c;
			16'hff44: y = 16'hff4d;
			16'hff45: y = 16'hff4d;
			16'hff46: y = 16'hff4e;
			16'hff47: y = 16'hff4f;
			16'hff48: y = 16'hff50;
			16'hff49: y = 16'hff51;
			16'hff4a: y = 16'hff52;
			16'hff4b: y = 16'hff53;
			16'hff4c: y = 16'hff54;
			16'hff4d: y = 16'hff54;
			16'hff4e: y = 16'hff55;
			16'hff4f: y = 16'hff56;
			16'hff50: y = 16'hff57;
			16'hff51: y = 16'hff58;
			16'hff52: y = 16'hff59;
			16'hff53: y = 16'hff5a;
			16'hff54: y = 16'hff5b;
			16'hff55: y = 16'hff5c;
			16'hff56: y = 16'hff5c;
			16'hff57: y = 16'hff5d;
			16'hff58: y = 16'hff5e;
			16'hff59: y = 16'hff5f;
			16'hff5a: y = 16'hff60;
			16'hff5b: y = 16'hff61;
			16'hff5c: y = 16'hff62;
			16'hff5d: y = 16'hff63;
			16'hff5e: y = 16'hff64;
			16'hff5f: y = 16'hff65;
			16'hff60: y = 16'hff66;
			16'hff61: y = 16'hff66;
			16'hff62: y = 16'hff67;
			16'hff63: y = 16'hff68;
			16'hff64: y = 16'hff69;
			16'hff65: y = 16'hff6a;
			16'hff66: y = 16'hff6b;
			16'hff67: y = 16'hff6c;
			16'hff68: y = 16'hff6d;
			16'hff69: y = 16'hff6e;
			16'hff6a: y = 16'hff6f;
			16'hff6b: y = 16'hff70;
			16'hff6c: y = 16'hff70;
			16'hff6d: y = 16'hff71;
			16'hff6e: y = 16'hff72;
			16'hff6f: y = 16'hff73;
			16'hff70: y = 16'hff74;
			16'hff71: y = 16'hff75;
			16'hff72: y = 16'hff76;
			16'hff73: y = 16'hff77;
			16'hff74: y = 16'hff78;
			16'hff75: y = 16'hff79;
			16'hff76: y = 16'hff7a;
			16'hff77: y = 16'hff7b;
			16'hff78: y = 16'hff7c;
			16'hff79: y = 16'hff7d;
			16'hff7a: y = 16'hff7d;
			16'hff7b: y = 16'hff7e;
			16'hff7c: y = 16'hff7f;
			16'hff7d: y = 16'hff80;
			16'hff7e: y = 16'hff81;
			16'hff7f: y = 16'hff82;
			16'hff80: y = 16'hff83;
			16'hff81: y = 16'hff84;
			16'hff82: y = 16'hff85;
			16'hff83: y = 16'hff86;
			16'hff84: y = 16'hff87;
			16'hff85: y = 16'hff88;
			16'hff86: y = 16'hff89;
			16'hff87: y = 16'hff8a;
			16'hff88: y = 16'hff8b;
			16'hff89: y = 16'hff8c;
			16'hff8a: y = 16'hff8d;
			16'hff8b: y = 16'hff8d;
			16'hff8c: y = 16'hff8e;
			16'hff8d: y = 16'hff8f;
			16'hff8e: y = 16'hff90;
			16'hff8f: y = 16'hff91;
			16'hff90: y = 16'hff92;
			16'hff91: y = 16'hff93;
			16'hff92: y = 16'hff94;
			16'hff93: y = 16'hff95;
			16'hff94: y = 16'hff96;
			16'hff95: y = 16'hff97;
			16'hff96: y = 16'hff98;
			16'hff97: y = 16'hff99;
			16'hff98: y = 16'hff9a;
			16'hff99: y = 16'hff9b;
			16'hff9a: y = 16'hff9c;
			16'hff9b: y = 16'hff9d;
			16'hff9c: y = 16'hff9e;
			16'hff9d: y = 16'hff9f;
			16'hff9e: y = 16'hffa0;
			16'hff9f: y = 16'hffa1;
			16'hffa0: y = 16'hffa2;
			16'hffa1: y = 16'hffa3;
			16'hffa2: y = 16'hffa4;
			16'hffa3: y = 16'hffa5;
			16'hffa4: y = 16'hffa5;
			16'hffa5: y = 16'hffa6;
			16'hffa6: y = 16'hffa7;
			16'hffa7: y = 16'hffa8;
			16'hffa8: y = 16'hffa9;
			16'hffa9: y = 16'hffaa;
			16'hffaa: y = 16'hffab;
			16'hffab: y = 16'hffac;
			16'hffac: y = 16'hffad;
			16'hffad: y = 16'hffae;
			16'hffae: y = 16'hffaf;
			16'hffaf: y = 16'hffb0;
			16'hffb0: y = 16'hffb1;
			16'hffb1: y = 16'hffb2;
			16'hffb2: y = 16'hffb3;
			16'hffb3: y = 16'hffb4;
			16'hffb4: y = 16'hffb5;
			16'hffb5: y = 16'hffb6;
			16'hffb6: y = 16'hffb7;
			16'hffb7: y = 16'hffb8;
			16'hffb8: y = 16'hffb9;
			16'hffb9: y = 16'hffba;
			16'hffba: y = 16'hffbb;
			16'hffbb: y = 16'hffbc;
			16'hffbc: y = 16'hffbd;
			16'hffbd: y = 16'hffbe;
			16'hffbe: y = 16'hffbf;
			16'hffbf: y = 16'hffc0;
			16'hffc0: y = 16'hffc1;
			16'hffc1: y = 16'hffc2;
			16'hffc2: y = 16'hffc3;
			16'hffc3: y = 16'hffc4;
			16'hffc4: y = 16'hffc5;
			16'hffc5: y = 16'hffc6;
			16'hffc6: y = 16'hffc7;
			16'hffc7: y = 16'hffc8;
			16'hffc8: y = 16'hffc9;
			16'hffc9: y = 16'hffca;
			16'hffca: y = 16'hffcb;
			16'hffcb: y = 16'hffcc;
			16'hffcc: y = 16'hffcd;
			16'hffcd: y = 16'hffce;
			16'hffce: y = 16'hffcf;
			16'hffcf: y = 16'hffd0;
			16'hffd0: y = 16'hffd1;
			16'hffd1: y = 16'hffd2;
			16'hffd2: y = 16'hffd3;
			16'hffd3: y = 16'hffd4;
			16'hffd4: y = 16'hffd5;
			16'hffd5: y = 16'hffd6;
			16'hffd6: y = 16'hffd7;
			16'hffd7: y = 16'hffd8;
			16'hffd8: y = 16'hffd9;
			16'hffd9: y = 16'hffda;
			16'hffda: y = 16'hffdb;
			16'hffdb: y = 16'hffdc;
			16'hffdc: y = 16'hffdd;
			16'hffdd: y = 16'hffde;
			16'hffde: y = 16'hffdf;
			16'hffdf: y = 16'hffe0;
			16'hffe0: y = 16'hffe1;
			16'hffe1: y = 16'hffe2;
			16'hffe2: y = 16'hffe3;
			16'hffe3: y = 16'hffe4;
			16'hffe4: y = 16'hffe5;
			16'hffe5: y = 16'hffe6;
			16'hffe6: y = 16'hffe7;
			16'hffe7: y = 16'hffe8;
			16'hffe8: y = 16'hffe9;
			16'hffe9: y = 16'hffea;
			16'hffea: y = 16'hffeb;
			16'hffeb: y = 16'hffec;
			16'hffec: y = 16'hffed;
			16'hffed: y = 16'hffee;
			16'hffee: y = 16'hffef;
			16'hffef: y = 16'hfff0;
			16'hfff0: y = 16'hfff1;
			16'hfff1: y = 16'hfff2;
			16'hfff2: y = 16'hfff3;
			16'hfff3: y = 16'hfff4;
			16'hfff4: y = 16'hfff5;
			16'hfff5: y = 16'hfff6;
			16'hfff6: y = 16'hfff7;
			16'hfff7: y = 16'hfff8;
			16'hfff8: y = 16'hfff9;
			16'hfff9: y = 16'hfffa;
			16'hfffa: y = 16'hfffb;
			16'hfffb: y = 16'hfffc;
			16'hfffc: y = 16'hfffd;
			16'hfffd: y = 16'hfffe;
			16'hfffe: y = 16'hffff;
			16'hffff: y = 16'h0;
			16'h0: y = 16'h0;
			16'h1: y = 16'h0;
			16'h2: y = 16'h1;
			16'h3: y = 16'h2;
			16'h4: y = 16'h3;
			16'h5: y = 16'h4;
			16'h6: y = 16'h5;
			16'h7: y = 16'h6;
			16'h8: y = 16'h7;
			16'h9: y = 16'h8;
			16'ha: y = 16'h9;
			16'hb: y = 16'ha;
			16'hc: y = 16'hb;
			16'hd: y = 16'hc;
			16'he: y = 16'hd;
			16'hf: y = 16'he;
			16'h10: y = 16'hf;
			16'h11: y = 16'h10;
			16'h12: y = 16'h11;
			16'h13: y = 16'h12;
			16'h14: y = 16'h13;
			16'h15: y = 16'h14;
			16'h16: y = 16'h15;
			16'h17: y = 16'h16;
			16'h18: y = 16'h17;
			16'h19: y = 16'h18;
			16'h1a: y = 16'h19;
			16'h1b: y = 16'h1a;
			16'h1c: y = 16'h1b;
			16'h1d: y = 16'h1c;
			16'h1e: y = 16'h1d;
			16'h1f: y = 16'h1e;
			16'h20: y = 16'h1f;
			16'h21: y = 16'h20;
			16'h22: y = 16'h21;
			16'h23: y = 16'h22;
			16'h24: y = 16'h23;
			16'h25: y = 16'h24;
			16'h26: y = 16'h25;
			16'h27: y = 16'h26;
			16'h28: y = 16'h27;
			16'h29: y = 16'h28;
			16'h2a: y = 16'h29;
			16'h2b: y = 16'h2a;
			16'h2c: y = 16'h2b;
			16'h2d: y = 16'h2c;
			16'h2e: y = 16'h2d;
			16'h2f: y = 16'h2e;
			16'h30: y = 16'h2f;
			16'h31: y = 16'h30;
			16'h32: y = 16'h31;
			16'h33: y = 16'h32;
			16'h34: y = 16'h33;
			16'h35: y = 16'h34;
			16'h36: y = 16'h35;
			16'h37: y = 16'h36;
			16'h38: y = 16'h37;
			16'h39: y = 16'h38;
			16'h3a: y = 16'h39;
			16'h3b: y = 16'h3a;
			16'h3c: y = 16'h3b;
			16'h3d: y = 16'h3c;
			16'h3e: y = 16'h3d;
			16'h3f: y = 16'h3e;
			16'h40: y = 16'h3f;
			16'h41: y = 16'h40;
			16'h42: y = 16'h41;
			16'h43: y = 16'h42;
			16'h44: y = 16'h43;
			16'h45: y = 16'h44;
			16'h46: y = 16'h45;
			16'h47: y = 16'h46;
			16'h48: y = 16'h47;
			16'h49: y = 16'h48;
			16'h4a: y = 16'h49;
			16'h4b: y = 16'h4a;
			16'h4c: y = 16'h4b;
			16'h4d: y = 16'h4c;
			16'h4e: y = 16'h4d;
			16'h4f: y = 16'h4e;
			16'h50: y = 16'h4f;
			16'h51: y = 16'h50;
			16'h52: y = 16'h51;
			16'h53: y = 16'h52;
			16'h54: y = 16'h53;
			16'h55: y = 16'h54;
			16'h56: y = 16'h55;
			16'h57: y = 16'h56;
			16'h58: y = 16'h57;
			16'h59: y = 16'h58;
			16'h5a: y = 16'h59;
			16'h5b: y = 16'h5a;
			16'h5c: y = 16'h5b;
			16'h5d: y = 16'h5b;
			16'h5e: y = 16'h5c;
			16'h5f: y = 16'h5d;
			16'h60: y = 16'h5e;
			16'h61: y = 16'h5f;
			16'h62: y = 16'h60;
			16'h63: y = 16'h61;
			16'h64: y = 16'h62;
			16'h65: y = 16'h63;
			16'h66: y = 16'h64;
			16'h67: y = 16'h65;
			16'h68: y = 16'h66;
			16'h69: y = 16'h67;
			16'h6a: y = 16'h68;
			16'h6b: y = 16'h69;
			16'h6c: y = 16'h6a;
			16'h6d: y = 16'h6b;
			16'h6e: y = 16'h6c;
			16'h6f: y = 16'h6d;
			16'h70: y = 16'h6e;
			16'h71: y = 16'h6f;
			16'h72: y = 16'h70;
			16'h73: y = 16'h71;
			16'h74: y = 16'h72;
			16'h75: y = 16'h73;
			16'h76: y = 16'h73;
			16'h77: y = 16'h74;
			16'h78: y = 16'h75;
			16'h79: y = 16'h76;
			16'h7a: y = 16'h77;
			16'h7b: y = 16'h78;
			16'h7c: y = 16'h79;
			16'h7d: y = 16'h7a;
			16'h7e: y = 16'h7b;
			16'h7f: y = 16'h7c;
			16'h80: y = 16'h7d;
			16'h81: y = 16'h7e;
			16'h82: y = 16'h7f;
			16'h83: y = 16'h80;
			16'h84: y = 16'h81;
			16'h85: y = 16'h82;
			16'h86: y = 16'h83;
			16'h87: y = 16'h83;
			16'h88: y = 16'h84;
			16'h89: y = 16'h85;
			16'h8a: y = 16'h86;
			16'h8b: y = 16'h87;
			16'h8c: y = 16'h88;
			16'h8d: y = 16'h89;
			16'h8e: y = 16'h8a;
			16'h8f: y = 16'h8b;
			16'h90: y = 16'h8c;
			16'h91: y = 16'h8d;
			16'h92: y = 16'h8e;
			16'h93: y = 16'h8f;
			16'h94: y = 16'h90;
			16'h95: y = 16'h90;
			16'h96: y = 16'h91;
			16'h97: y = 16'h92;
			16'h98: y = 16'h93;
			16'h99: y = 16'h94;
			16'h9a: y = 16'h95;
			16'h9b: y = 16'h96;
			16'h9c: y = 16'h97;
			16'h9d: y = 16'h98;
			16'h9e: y = 16'h99;
			16'h9f: y = 16'h9a;
			16'ha0: y = 16'h9a;
			16'ha1: y = 16'h9b;
			16'ha2: y = 16'h9c;
			16'ha3: y = 16'h9d;
			16'ha4: y = 16'h9e;
			16'ha5: y = 16'h9f;
			16'ha6: y = 16'ha0;
			16'ha7: y = 16'ha1;
			16'ha8: y = 16'ha2;
			16'ha9: y = 16'ha3;
			16'haa: y = 16'ha4;
			16'hab: y = 16'ha4;
			16'hac: y = 16'ha5;
			16'had: y = 16'ha6;
			16'hae: y = 16'ha7;
			16'haf: y = 16'ha8;
			16'hb0: y = 16'ha9;
			16'hb1: y = 16'haa;
			16'hb2: y = 16'hab;
			16'hb3: y = 16'hac;
			16'hb4: y = 16'hac;
			16'hb5: y = 16'had;
			16'hb6: y = 16'hae;
			16'hb7: y = 16'haf;
			16'hb8: y = 16'hb0;
			16'hb9: y = 16'hb1;
			16'hba: y = 16'hb2;
			16'hbb: y = 16'hb3;
			16'hbc: y = 16'hb3;
			16'hbd: y = 16'hb4;
			16'hbe: y = 16'hb5;
			16'hbf: y = 16'hb6;
			16'hc0: y = 16'hb7;
			16'hc1: y = 16'hb8;
			16'hc2: y = 16'hb9;
			16'hc3: y = 16'hba;
			16'hc4: y = 16'hba;
			16'hc5: y = 16'hbb;
			16'hc6: y = 16'hbc;
			16'hc7: y = 16'hbd;
			16'hc8: y = 16'hbe;
			16'hc9: y = 16'hbf;
			16'hca: y = 16'hc0;
			16'hcb: y = 16'hc0;
			16'hcc: y = 16'hc1;
			16'hcd: y = 16'hc2;
			16'hce: y = 16'hc3;
			16'hcf: y = 16'hc4;
			16'hd0: y = 16'hc5;
			16'hd1: y = 16'hc6;
			16'hd2: y = 16'hc6;
			16'hd3: y = 16'hc7;
			16'hd4: y = 16'hc8;
			16'hd5: y = 16'hc9;
			16'hd6: y = 16'hca;
			16'hd7: y = 16'hcb;
			16'hd8: y = 16'hcc;
			16'hd9: y = 16'hcc;
			16'hda: y = 16'hcd;
			16'hdb: y = 16'hce;
			16'hdc: y = 16'hcf;
			16'hdd: y = 16'hd0;
			16'hde: y = 16'hd1;
			16'hdf: y = 16'hd1;
			16'he0: y = 16'hd2;
			16'he1: y = 16'hd3;
			16'he2: y = 16'hd4;
			16'he3: y = 16'hd5;
			16'he4: y = 16'hd6;
			16'he5: y = 16'hd6;
			16'he6: y = 16'hd7;
			16'he7: y = 16'hd8;
			16'he8: y = 16'hd9;
			16'he9: y = 16'hda;
			16'hea: y = 16'hda;
			16'heb: y = 16'hdb;
			16'hec: y = 16'hdc;
			16'hed: y = 16'hdd;
			16'hee: y = 16'hde;
			16'hef: y = 16'hdf;
			16'hf0: y = 16'hdf;
			16'hf1: y = 16'he0;
			16'hf2: y = 16'he1;
			16'hf3: y = 16'he2;
			16'hf4: y = 16'he3;
			16'hf5: y = 16'he3;
			16'hf6: y = 16'he4;
			16'hf7: y = 16'he5;
			16'hf8: y = 16'he6;
			16'hf9: y = 16'he7;
			16'hfa: y = 16'he7;
			16'hfb: y = 16'he8;
			16'hfc: y = 16'he9;
			16'hfd: y = 16'hea;
			16'hfe: y = 16'heb;
			16'hff: y = 16'heb;
			16'h100: y = 16'hec;
			16'h101: y = 16'hed;
			16'h102: y = 16'hee;
			16'h103: y = 16'hee;
			16'h104: y = 16'hef;
			16'h105: y = 16'hf0;
			16'h106: y = 16'hf1;
			16'h107: y = 16'hf2;
			16'h108: y = 16'hf2;
			16'h109: y = 16'hf3;
			16'h10a: y = 16'hf4;
			16'h10b: y = 16'hf5;
			16'h10c: y = 16'hf5;
			16'h10d: y = 16'hf6;
			16'h10e: y = 16'hf7;
			16'h10f: y = 16'hf8;
			16'h110: y = 16'hf9;
			16'h111: y = 16'hf9;
			16'h112: y = 16'hfa;
			16'h113: y = 16'hfb;
			16'h114: y = 16'hfc;
			16'h115: y = 16'hfc;
			16'h116: y = 16'hfd;
			16'h117: y = 16'hfe;
			16'h118: y = 16'hff;
			16'h119: y = 16'hff;
			16'h11a: y = 16'h100;
			16'h11b: y = 16'h101;
			16'h11c: y = 16'h102;
			16'h11d: y = 16'h102;
			16'h11e: y = 16'h103;
			16'h11f: y = 16'h104;
			16'h120: y = 16'h105;
			16'h121: y = 16'h105;
			16'h122: y = 16'h106;
			16'h123: y = 16'h107;
			16'h124: y = 16'h107;
			16'h125: y = 16'h108;
			16'h126: y = 16'h109;
			16'h127: y = 16'h10a;
			16'h128: y = 16'h10a;
			16'h129: y = 16'h10b;
			16'h12a: y = 16'h10c;
			16'h12b: y = 16'h10d;
			16'h12c: y = 16'h10d;
			16'h12d: y = 16'h10e;
			16'h12e: y = 16'h10f;
			16'h12f: y = 16'h10f;
			16'h130: y = 16'h110;
			16'h131: y = 16'h111;
			16'h132: y = 16'h112;
			16'h133: y = 16'h112;
			16'h134: y = 16'h113;
			16'h135: y = 16'h114;
			16'h136: y = 16'h114;
			16'h137: y = 16'h115;
			16'h138: y = 16'h116;
			16'h139: y = 16'h117;
			16'h13a: y = 16'h117;
			16'h13b: y = 16'h118;
			16'h13c: y = 16'h119;
			16'h13d: y = 16'h119;
			16'h13e: y = 16'h11a;
			16'h13f: y = 16'h11b;
			16'h140: y = 16'h11b;
			16'h141: y = 16'h11c;
			16'h142: y = 16'h11d;
			16'h143: y = 16'h11e;
			16'h144: y = 16'h11e;
			16'h145: y = 16'h11f;
			16'h146: y = 16'h120;
			16'h147: y = 16'h120;
			16'h148: y = 16'h121;
			16'h149: y = 16'h122;
			16'h14a: y = 16'h122;
			16'h14b: y = 16'h123;
			16'h14c: y = 16'h124;
			16'h14d: y = 16'h124;
			16'h14e: y = 16'h125;
			16'h14f: y = 16'h126;
			16'h150: y = 16'h126;
			16'h151: y = 16'h127;
			16'h152: y = 16'h128;
			16'h153: y = 16'h128;
			16'h154: y = 16'h129;
			16'h155: y = 16'h12a;
			16'h156: y = 16'h12a;
			16'h157: y = 16'h12b;
			16'h158: y = 16'h12c;
			16'h159: y = 16'h12c;
			16'h15a: y = 16'h12d;
			16'h15b: y = 16'h12e;
			16'h15c: y = 16'h12e;
			16'h15d: y = 16'h12f;
			16'h15e: y = 16'h130;
			16'h15f: y = 16'h130;
			16'h160: y = 16'h131;
			16'h161: y = 16'h131;
			16'h162: y = 16'h132;
			16'h163: y = 16'h133;
			16'h164: y = 16'h133;
			16'h165: y = 16'h134;
			16'h166: y = 16'h135;
			16'h167: y = 16'h135;
			16'h168: y = 16'h136;
			16'h169: y = 16'h137;
			16'h16a: y = 16'h137;
			16'h16b: y = 16'h138;
			16'h16c: y = 16'h138;
			16'h16d: y = 16'h139;
			16'h16e: y = 16'h13a;
			16'h16f: y = 16'h13a;
			16'h170: y = 16'h13b;
			16'h171: y = 16'h13c;
			16'h172: y = 16'h13c;
			16'h173: y = 16'h13d;
			16'h174: y = 16'h13d;
			16'h175: y = 16'h13e;
			16'h176: y = 16'h13f;
			16'h177: y = 16'h13f;
			16'h178: y = 16'h140;
			16'h179: y = 16'h140;
			16'h17a: y = 16'h141;
			16'h17b: y = 16'h142;
			16'h17c: y = 16'h142;
			16'h17d: y = 16'h143;
			16'h17e: y = 16'h144;
			16'h17f: y = 16'h144;
			16'h180: y = 16'h145;
			16'h181: y = 16'h145;
			16'h182: y = 16'h146;
			16'h183: y = 16'h146;
			16'h184: y = 16'h147;
			16'h185: y = 16'h148;
			16'h186: y = 16'h148;
			16'h187: y = 16'h149;
			16'h188: y = 16'h149;
			16'h189: y = 16'h14a;
			16'h18a: y = 16'h14b;
			16'h18b: y = 16'h14b;
			16'h18c: y = 16'h14c;
			16'h18d: y = 16'h14c;
			16'h18e: y = 16'h14d;
			16'h18f: y = 16'h14d;
			16'h190: y = 16'h14e;
			16'h191: y = 16'h14f;
			16'h192: y = 16'h14f;
			16'h193: y = 16'h150;
			16'h194: y = 16'h150;
			16'h195: y = 16'h151;
			16'h196: y = 16'h151;
			16'h197: y = 16'h152;
			16'h198: y = 16'h153;
			16'h199: y = 16'h153;
			16'h19a: y = 16'h154;
			16'h19b: y = 16'h154;
			16'h19c: y = 16'h155;
			16'h19d: y = 16'h155;
			16'h19e: y = 16'h156;
			16'h19f: y = 16'h156;
			16'h1a0: y = 16'h157;
			16'h1a1: y = 16'h158;
			16'h1a2: y = 16'h158;
			16'h1a3: y = 16'h159;
			16'h1a4: y = 16'h159;
			16'h1a5: y = 16'h15a;
			16'h1a6: y = 16'h15a;
			16'h1a7: y = 16'h15b;
			16'h1a8: y = 16'h15b;
			16'h1a9: y = 16'h15c;
			16'h1aa: y = 16'h15c;
			16'h1ab: y = 16'h15d;
			16'h1ac: y = 16'h15e;
			16'h1ad: y = 16'h15e;
			16'h1ae: y = 16'h15f;
			16'h1af: y = 16'h15f;
			16'h1b0: y = 16'h160;
			16'h1b1: y = 16'h160;
			16'h1b2: y = 16'h161;
			16'h1b3: y = 16'h161;
			16'h1b4: y = 16'h162;
			16'h1b5: y = 16'h162;
			16'h1b6: y = 16'h163;
			16'h1b7: y = 16'h163;
			16'h1b8: y = 16'h164;
			16'h1b9: y = 16'h164;
			16'h1ba: y = 16'h165;
			16'h1bb: y = 16'h165;
			16'h1bc: y = 16'h166;
			16'h1bd: y = 16'h166;
			16'h1be: y = 16'h167;
			16'h1bf: y = 16'h167;
			16'h1c0: y = 16'h168;
			16'h1c1: y = 16'h168;
			16'h1c2: y = 16'h169;
			16'h1c3: y = 16'h169;
			16'h1c4: y = 16'h16a;
			16'h1c5: y = 16'h16a;
			16'h1c6: y = 16'h16b;
			16'h1c7: y = 16'h16b;
			16'h1c8: y = 16'h16c;
			16'h1c9: y = 16'h16c;
			16'h1ca: y = 16'h16d;
			16'h1cb: y = 16'h16d;
			16'h1cc: y = 16'h16e;
			16'h1cd: y = 16'h16e;
			16'h1ce: y = 16'h16f;
			16'h1cf: y = 16'h16f;
			16'h1d0: y = 16'h170;
			16'h1d1: y = 16'h170;
			16'h1d2: y = 16'h171;
			16'h1d3: y = 16'h171;
			16'h1d4: y = 16'h172;
			16'h1d5: y = 16'h172;
			16'h1d6: y = 16'h173;
			16'h1d7: y = 16'h173;
			16'h1d8: y = 16'h174;
			16'h1d9: y = 16'h174;
			16'h1da: y = 16'h175;
			16'h1db: y = 16'h175;
			16'h1dc: y = 16'h175;
			16'h1dd: y = 16'h176;
			16'h1de: y = 16'h176;
			16'h1df: y = 16'h177;
			16'h1e0: y = 16'h177;
			16'h1e1: y = 16'h178;
			16'h1e2: y = 16'h178;
			16'h1e3: y = 16'h179;
			16'h1e4: y = 16'h179;
			16'h1e5: y = 16'h17a;
			16'h1e6: y = 16'h17a;
			16'h1e7: y = 16'h17b;
			16'h1e8: y = 16'h17b;
			16'h1e9: y = 16'h17b;
			16'h1ea: y = 16'h17c;
			16'h1eb: y = 16'h17c;
			16'h1ec: y = 16'h17d;
			16'h1ed: y = 16'h17d;
			16'h1ee: y = 16'h17e;
			16'h1ef: y = 16'h17e;
			16'h1f0: y = 16'h17f;
			16'h1f1: y = 16'h17f;
			16'h1f2: y = 16'h17f;
			16'h1f3: y = 16'h180;
			16'h1f4: y = 16'h180;
			16'h1f5: y = 16'h181;
			16'h1f6: y = 16'h181;
			16'h1f7: y = 16'h182;
			16'h1f8: y = 16'h182;
			16'h1f9: y = 16'h182;
			16'h1fa: y = 16'h183;
			16'h1fb: y = 16'h183;
			16'h1fc: y = 16'h184;
			16'h1fd: y = 16'h184;
			16'h1fe: y = 16'h185;
			16'h1ff: y = 16'h185;
			16'h200: y = 16'h185;
			16'h201: y = 16'h186;
			16'h202: y = 16'h186;
			16'h203: y = 16'h187;
			16'h204: y = 16'h187;
			16'h205: y = 16'h188;
			16'h206: y = 16'h188;
			16'h207: y = 16'h188;
			16'h208: y = 16'h189;
			16'h209: y = 16'h189;
			16'h20a: y = 16'h18a;
			16'h20b: y = 16'h18a;
			16'h20c: y = 16'h18a;
			16'h20d: y = 16'h18b;
			16'h20e: y = 16'h18b;
			16'h20f: y = 16'h18c;
			16'h210: y = 16'h18c;
			16'h211: y = 16'h18c;
			16'h212: y = 16'h18d;
			16'h213: y = 16'h18d;
			16'h214: y = 16'h18e;
			16'h215: y = 16'h18e;
			16'h216: y = 16'h18e;
			16'h217: y = 16'h18f;
			16'h218: y = 16'h18f;
			16'h219: y = 16'h190;
			16'h21a: y = 16'h190;
			16'h21b: y = 16'h190;
			16'h21c: y = 16'h191;
			16'h21d: y = 16'h191;
			16'h21e: y = 16'h191;
			16'h21f: y = 16'h192;
			16'h220: y = 16'h192;
			16'h221: y = 16'h193;
			16'h222: y = 16'h193;
			16'h223: y = 16'h193;
			16'h224: y = 16'h194;
			16'h225: y = 16'h194;
			16'h226: y = 16'h195;
			16'h227: y = 16'h195;
			16'h228: y = 16'h195;
			16'h229: y = 16'h196;
			16'h22a: y = 16'h196;
			16'h22b: y = 16'h196;
			16'h22c: y = 16'h197;
			16'h22d: y = 16'h197;
			16'h22e: y = 16'h197;
			16'h22f: y = 16'h198;
			16'h230: y = 16'h198;
			16'h231: y = 16'h199;
			16'h232: y = 16'h199;
			16'h233: y = 16'h199;
			16'h234: y = 16'h19a;
			16'h235: y = 16'h19a;
			16'h236: y = 16'h19a;
			16'h237: y = 16'h19b;
			16'h238: y = 16'h19b;
			16'h239: y = 16'h19b;
			16'h23a: y = 16'h19c;
			16'h23b: y = 16'h19c;
			16'h23c: y = 16'h19c;
			16'h23d: y = 16'h19d;
			16'h23e: y = 16'h19d;
			16'h23f: y = 16'h19e;
			16'h240: y = 16'h19e;
			16'h241: y = 16'h19e;
			16'h242: y = 16'h19f;
			16'h243: y = 16'h19f;
			16'h244: y = 16'h19f;
			16'h245: y = 16'h1a0;
			16'h246: y = 16'h1a0;
			16'h247: y = 16'h1a0;
			16'h248: y = 16'h1a1;
			16'h249: y = 16'h1a1;
			16'h24a: y = 16'h1a1;
			16'h24b: y = 16'h1a2;
			16'h24c: y = 16'h1a2;
			16'h24d: y = 16'h1a2;
			16'h24e: y = 16'h1a3;
			16'h24f: y = 16'h1a3;
			16'h250: y = 16'h1a3;
			16'h251: y = 16'h1a4;
			16'h252: y = 16'h1a4;
			16'h253: y = 16'h1a4;
			16'h254: y = 16'h1a5;
			16'h255: y = 16'h1a5;
			16'h256: y = 16'h1a5;
			16'h257: y = 16'h1a6;
			16'h258: y = 16'h1a6;
			16'h259: y = 16'h1a6;
			16'h25a: y = 16'h1a6;
			16'h25b: y = 16'h1a7;
			16'h25c: y = 16'h1a7;
			16'h25d: y = 16'h1a7;
			16'h25e: y = 16'h1a8;
			16'h25f: y = 16'h1a8;
			16'h260: y = 16'h1a8;
			16'h261: y = 16'h1a9;
			16'h262: y = 16'h1a9;
			16'h263: y = 16'h1a9;
			16'h264: y = 16'h1aa;
			16'h265: y = 16'h1aa;
			16'h266: y = 16'h1aa;
			16'h267: y = 16'h1ab;
			16'h268: y = 16'h1ab;
			16'h269: y = 16'h1ab;
			16'h26a: y = 16'h1ab;
			16'h26b: y = 16'h1ac;
			16'h26c: y = 16'h1ac;
			16'h26d: y = 16'h1ac;
			16'h26e: y = 16'h1ad;
			16'h26f: y = 16'h1ad;
			16'h270: y = 16'h1ad;
			16'h271: y = 16'h1ae;
			16'h272: y = 16'h1ae;
			16'h273: y = 16'h1ae;
			16'h274: y = 16'h1ae;
			16'h275: y = 16'h1af;
			16'h276: y = 16'h1af;
			16'h277: y = 16'h1af;
			16'h278: y = 16'h1b0;
			16'h279: y = 16'h1b0;
			16'h27a: y = 16'h1b0;
			16'h27b: y = 16'h1b0;
			16'h27c: y = 16'h1b1;
			16'h27d: y = 16'h1b1;
			16'h27e: y = 16'h1b1;
			16'h27f: y = 16'h1b2;
			16'h280: y = 16'h1b2;
			16'h281: y = 16'h1b2;
			16'h282: y = 16'h1b2;
			16'h283: y = 16'h1b3;
			16'h284: y = 16'h1b3;
			16'h285: y = 16'h1b3;
			16'h286: y = 16'h1b3;
			16'h287: y = 16'h1b4;
			16'h288: y = 16'h1b4;
			16'h289: y = 16'h1b4;
			16'h28a: y = 16'h1b5;
			16'h28b: y = 16'h1b5;
			16'h28c: y = 16'h1b5;
			16'h28d: y = 16'h1b5;
			16'h28e: y = 16'h1b6;
			16'h28f: y = 16'h1b6;
			16'h290: y = 16'h1b6;
			16'h291: y = 16'h1b6;
			16'h292: y = 16'h1b7;
			16'h293: y = 16'h1b7;
			16'h294: y = 16'h1b7;
			16'h295: y = 16'h1b8;
			16'h296: y = 16'h1b8;
			16'h297: y = 16'h1b8;
			16'h298: y = 16'h1b8;
			16'h299: y = 16'h1b9;
			16'h29a: y = 16'h1b9;
			16'h29b: y = 16'h1b9;
			16'h29c: y = 16'h1b9;
			16'h29d: y = 16'h1ba;
			16'h29e: y = 16'h1ba;
			16'h29f: y = 16'h1ba;
			16'h2a0: y = 16'h1ba;
			16'h2a1: y = 16'h1bb;
			16'h2a2: y = 16'h1bb;
			16'h2a3: y = 16'h1bb;
			16'h2a4: y = 16'h1bb;
			16'h2a5: y = 16'h1bc;
			16'h2a6: y = 16'h1bc;
			16'h2a7: y = 16'h1bc;
			16'h2a8: y = 16'h1bc;
			16'h2a9: y = 16'h1bd;
			16'h2aa: y = 16'h1bd;
			16'h2ab: y = 16'h1bd;
			16'h2ac: y = 16'h1bd;
			16'h2ad: y = 16'h1be;
			16'h2ae: y = 16'h1be;
			16'h2af: y = 16'h1be;
			16'h2b0: y = 16'h1be;
			16'h2b1: y = 16'h1be;
			16'h2b2: y = 16'h1bf;
			16'h2b3: y = 16'h1bf;
			16'h2b4: y = 16'h1bf;
			16'h2b5: y = 16'h1bf;
			16'h2b6: y = 16'h1c0;
			16'h2b7: y = 16'h1c0;
			16'h2b8: y = 16'h1c0;
			16'h2b9: y = 16'h1c0;
			16'h2ba: y = 16'h1c1;
			16'h2bb: y = 16'h1c1;
			16'h2bc: y = 16'h1c1;
			16'h2bd: y = 16'h1c1;
			16'h2be: y = 16'h1c2;
			16'h2bf: y = 16'h1c2;
			16'h2c0: y = 16'h1c2;
			16'h2c1: y = 16'h1c2;
			16'h2c2: y = 16'h1c2;
			16'h2c3: y = 16'h1c3;
			16'h2c4: y = 16'h1c3;
			16'h2c5: y = 16'h1c3;
			16'h2c6: y = 16'h1c3;
			16'h2c7: y = 16'h1c4;
			16'h2c8: y = 16'h1c4;
			16'h2c9: y = 16'h1c4;
			16'h2ca: y = 16'h1c4;
			16'h2cb: y = 16'h1c4;
			16'h2cc: y = 16'h1c5;
			16'h2cd: y = 16'h1c5;
			16'h2ce: y = 16'h1c5;
			16'h2cf: y = 16'h1c5;
			16'h2d0: y = 16'h1c5;
			16'h2d1: y = 16'h1c6;
			16'h2d2: y = 16'h1c6;
			16'h2d3: y = 16'h1c6;
			16'h2d4: y = 16'h1c6;
			16'h2d5: y = 16'h1c7;
			16'h2d6: y = 16'h1c7;
			16'h2d7: y = 16'h1c7;
			16'h2d8: y = 16'h1c7;
			16'h2d9: y = 16'h1c7;
			16'h2da: y = 16'h1c8;
			16'h2db: y = 16'h1c8;
			16'h2dc: y = 16'h1c8;
			16'h2dd: y = 16'h1c8;
			16'h2de: y = 16'h1c8;
			16'h2df: y = 16'h1c9;
			16'h2e0: y = 16'h1c9;
			16'h2e1: y = 16'h1c9;
			16'h2e2: y = 16'h1c9;
			16'h2e3: y = 16'h1c9;
			16'h2e4: y = 16'h1ca;
			16'h2e5: y = 16'h1ca;
			16'h2e6: y = 16'h1ca;
			16'h2e7: y = 16'h1ca;
			16'h2e8: y = 16'h1ca;
			16'h2e9: y = 16'h1cb;
			16'h2ea: y = 16'h1cb;
			16'h2eb: y = 16'h1cb;
			16'h2ec: y = 16'h1cb;
			16'h2ed: y = 16'h1cb;
			16'h2ee: y = 16'h1cc;
			16'h2ef: y = 16'h1cc;
			16'h2f0: y = 16'h1cc;
			16'h2f1: y = 16'h1cc;
			16'h2f2: y = 16'h1cc;
			16'h2f3: y = 16'h1cd;
			16'h2f4: y = 16'h1cd;
			16'h2f5: y = 16'h1cd;
			16'h2f6: y = 16'h1cd;
			16'h2f7: y = 16'h1cd;
			16'h2f8: y = 16'h1cd;
			16'h2f9: y = 16'h1ce;
			16'h2fa: y = 16'h1ce;
			16'h2fb: y = 16'h1ce;
			16'h2fc: y = 16'h1ce;
			16'h2fd: y = 16'h1ce;
			16'h2fe: y = 16'h1cf;
			16'h2ff: y = 16'h1cf;
			16'h300: y = 16'h1cf;
			16'h301: y = 16'h1cf;
			16'h302: y = 16'h1cf;
			16'h303: y = 16'h1cf;
			16'h304: y = 16'h1d0;
			16'h305: y = 16'h1d0;
			16'h306: y = 16'h1d0;
			16'h307: y = 16'h1d0;
			16'h308: y = 16'h1d0;
			16'h309: y = 16'h1d1;
			16'h30a: y = 16'h1d1;
			16'h30b: y = 16'h1d1;
			16'h30c: y = 16'h1d1;
			16'h30d: y = 16'h1d1;
			16'h30e: y = 16'h1d1;
			16'h30f: y = 16'h1d2;
			16'h310: y = 16'h1d2;
			16'h311: y = 16'h1d2;
			16'h312: y = 16'h1d2;
			16'h313: y = 16'h1d2;
			16'h314: y = 16'h1d2;
			16'h315: y = 16'h1d3;
			16'h316: y = 16'h1d3;
			16'h317: y = 16'h1d3;
			16'h318: y = 16'h1d3;
			16'h319: y = 16'h1d3;
			16'h31a: y = 16'h1d3;
			16'h31b: y = 16'h1d4;
			16'h31c: y = 16'h1d4;
			16'h31d: y = 16'h1d4;
			16'h31e: y = 16'h1d4;
			16'h31f: y = 16'h1d4;
			16'h320: y = 16'h1d4;
			16'h321: y = 16'h1d5;
			16'h322: y = 16'h1d5;
			16'h323: y = 16'h1d5;
			16'h324: y = 16'h1d5;
			16'h325: y = 16'h1d5;
			16'h326: y = 16'h1d5;
			16'h327: y = 16'h1d6;
			16'h328: y = 16'h1d6;
			16'h329: y = 16'h1d6;
			16'h32a: y = 16'h1d6;
			16'h32b: y = 16'h1d6;
			16'h32c: y = 16'h1d6;
			16'h32d: y = 16'h1d6;
			16'h32e: y = 16'h1d7;
			16'h32f: y = 16'h1d7;
			16'h330: y = 16'h1d7;
			16'h331: y = 16'h1d7;
			16'h332: y = 16'h1d7;
			16'h333: y = 16'h1d7;
			16'h334: y = 16'h1d8;
			16'h335: y = 16'h1d8;
			16'h336: y = 16'h1d8;
			16'h337: y = 16'h1d8;
			16'h338: y = 16'h1d8;
			16'h339: y = 16'h1d8;
			16'h33a: y = 16'h1d8;
			16'h33b: y = 16'h1d9;
			16'h33c: y = 16'h1d9;
			16'h33d: y = 16'h1d9;
			16'h33e: y = 16'h1d9;
			16'h33f: y = 16'h1d9;
			16'h340: y = 16'h1d9;
			16'h341: y = 16'h1d9;
			16'h342: y = 16'h1da;
			16'h343: y = 16'h1da;
			16'h344: y = 16'h1da;
			16'h345: y = 16'h1da;
			16'h346: y = 16'h1da;
			16'h347: y = 16'h1da;
			16'h348: y = 16'h1da;
			16'h349: y = 16'h1db;
			16'h34a: y = 16'h1db;
			16'h34b: y = 16'h1db;
			16'h34c: y = 16'h1db;
			16'h34d: y = 16'h1db;
			16'h34e: y = 16'h1db;
			16'h34f: y = 16'h1db;
			16'h350: y = 16'h1dc;
			16'h351: y = 16'h1dc;
			16'h352: y = 16'h1dc;
			16'h353: y = 16'h1dc;
			16'h354: y = 16'h1dc;
			16'h355: y = 16'h1dc;
			16'h356: y = 16'h1dc;
			16'h357: y = 16'h1dc;
			16'h358: y = 16'h1dd;
			16'h359: y = 16'h1dd;
			16'h35a: y = 16'h1dd;
			16'h35b: y = 16'h1dd;
			16'h35c: y = 16'h1dd;
			16'h35d: y = 16'h1dd;
			16'h35e: y = 16'h1dd;
			16'h35f: y = 16'h1dd;
			16'h360: y = 16'h1de;
			16'h361: y = 16'h1de;
			16'h362: y = 16'h1de;
			16'h363: y = 16'h1de;
			16'h364: y = 16'h1de;
			16'h365: y = 16'h1de;
			16'h366: y = 16'h1de;
			16'h367: y = 16'h1df;
			16'h368: y = 16'h1df;
			16'h369: y = 16'h1df;
			16'h36a: y = 16'h1df;
			16'h36b: y = 16'h1df;
			16'h36c: y = 16'h1df;
			16'h36d: y = 16'h1df;
			16'h36e: y = 16'h1df;
			16'h36f: y = 16'h1df;
			16'h370: y = 16'h1e0;
			16'h371: y = 16'h1e0;
			16'h372: y = 16'h1e0;
			16'h373: y = 16'h1e0;
			16'h374: y = 16'h1e0;
			16'h375: y = 16'h1e0;
			16'h376: y = 16'h1e0;
			16'h377: y = 16'h1e0;
			16'h378: y = 16'h1e1;
			16'h379: y = 16'h1e1;
			16'h37a: y = 16'h1e1;
			16'h37b: y = 16'h1e1;
			16'h37c: y = 16'h1e1;
			16'h37d: y = 16'h1e1;
			16'h37e: y = 16'h1e1;
			16'h37f: y = 16'h1e1;
			16'h380: y = 16'h1e1;
			16'h381: y = 16'h1e2;
			16'h382: y = 16'h1e2;
			16'h383: y = 16'h1e2;
			16'h384: y = 16'h1e2;
			16'h385: y = 16'h1e2;
			16'h386: y = 16'h1e2;
			16'h387: y = 16'h1e2;
			16'h388: y = 16'h1e2;
			16'h389: y = 16'h1e2;
			16'h38a: y = 16'h1e3;
			16'h38b: y = 16'h1e3;
			16'h38c: y = 16'h1e3;
			16'h38d: y = 16'h1e3;
			16'h38e: y = 16'h1e3;
			16'h38f: y = 16'h1e3;
			16'h390: y = 16'h1e3;
			16'h391: y = 16'h1e3;
			16'h392: y = 16'h1e3;
			16'h393: y = 16'h1e4;
			16'h394: y = 16'h1e4;
			16'h395: y = 16'h1e4;
			16'h396: y = 16'h1e4;
			16'h397: y = 16'h1e4;
			16'h398: y = 16'h1e4;
			16'h399: y = 16'h1e4;
			16'h39a: y = 16'h1e4;
			16'h39b: y = 16'h1e4;
			16'h39c: y = 16'h1e5;
			16'h39d: y = 16'h1e5;
			16'h39e: y = 16'h1e5;
			16'h39f: y = 16'h1e5;
			16'h3a0: y = 16'h1e5;
			16'h3a1: y = 16'h1e5;
			16'h3a2: y = 16'h1e5;
			16'h3a3: y = 16'h1e5;
			16'h3a4: y = 16'h1e5;
			16'h3a5: y = 16'h1e5;
			16'h3a6: y = 16'h1e6;
			16'h3a7: y = 16'h1e6;
			16'h3a8: y = 16'h1e6;
			16'h3a9: y = 16'h1e6;
			16'h3aa: y = 16'h1e6;
			16'h3ab: y = 16'h1e6;
			16'h3ac: y = 16'h1e6;
			16'h3ad: y = 16'h1e6;
			16'h3ae: y = 16'h1e6;
			16'h3af: y = 16'h1e6;
			16'h3b0: y = 16'h1e6;
			16'h3b1: y = 16'h1e7;
			16'h3b2: y = 16'h1e7;
			16'h3b3: y = 16'h1e7;
			16'h3b4: y = 16'h1e7;
			16'h3b5: y = 16'h1e7;
			16'h3b6: y = 16'h1e7;
			16'h3b7: y = 16'h1e7;
			16'h3b8: y = 16'h1e7;
			16'h3b9: y = 16'h1e7;
			16'h3ba: y = 16'h1e7;
			16'h3bb: y = 16'h1e8;
			16'h3bc: y = 16'h1e8;
			16'h3bd: y = 16'h1e8;
			16'h3be: y = 16'h1e8;
			16'h3bf: y = 16'h1e8;
			16'h3c0: y = 16'h1e8;
			16'h3c1: y = 16'h1e8;
			16'h3c2: y = 16'h1e8;
			16'h3c3: y = 16'h1e8;
			16'h3c4: y = 16'h1e8;
			16'h3c5: y = 16'h1e8;
			16'h3c6: y = 16'h1e9;
			16'h3c7: y = 16'h1e9;
			16'h3c8: y = 16'h1e9;
			16'h3c9: y = 16'h1e9;
			16'h3ca: y = 16'h1e9;
			16'h3cb: y = 16'h1e9;
			16'h3cc: y = 16'h1e9;
			16'h3cd: y = 16'h1e9;
			16'h3ce: y = 16'h1e9;
			16'h3cf: y = 16'h1e9;
			16'h3d0: y = 16'h1e9;
			16'h3d1: y = 16'h1e9;
			16'h3d2: y = 16'h1ea;
			16'h3d3: y = 16'h1ea;
			16'h3d4: y = 16'h1ea;
			16'h3d5: y = 16'h1ea;
			16'h3d6: y = 16'h1ea;
			16'h3d7: y = 16'h1ea;
			16'h3d8: y = 16'h1ea;
			16'h3d9: y = 16'h1ea;
			16'h3da: y = 16'h1ea;
			16'h3db: y = 16'h1ea;
			16'h3dc: y = 16'h1ea;
			16'h3dd: y = 16'h1ea;
			16'h3de: y = 16'h1eb;
			16'h3df: y = 16'h1eb;
			16'h3e0: y = 16'h1eb;
			16'h3e1: y = 16'h1eb;
			16'h3e2: y = 16'h1eb;
			16'h3e3: y = 16'h1eb;
			16'h3e4: y = 16'h1eb;
			16'h3e5: y = 16'h1eb;
			16'h3e6: y = 16'h1eb;
			16'h3e7: y = 16'h1eb;
			16'h3e8: y = 16'h1eb;
			16'h3e9: y = 16'h1eb;
			16'h3ea: y = 16'h1eb;
			16'h3eb: y = 16'h1ec;
			16'h3ec: y = 16'h1ec;
			16'h3ed: y = 16'h1ec;
			16'h3ee: y = 16'h1ec;
			16'h3ef: y = 16'h1ec;
			16'h3f0: y = 16'h1ec;
			16'h3f1: y = 16'h1ec;
			16'h3f2: y = 16'h1ec;
			16'h3f3: y = 16'h1ec;
			16'h3f4: y = 16'h1ec;
			16'h3f5: y = 16'h1ec;
			16'h3f6: y = 16'h1ec;
			16'h3f7: y = 16'h1ec;
			16'h3f8: y = 16'h1ed;
			16'h3f9: y = 16'h1ed;
			16'h3fa: y = 16'h1ed;
			16'h3fb: y = 16'h1ed;
			16'h3fc: y = 16'h1ed;
			16'h3fd: y = 16'h1ed;
			16'h3fe: y = 16'h1ed;
			16'h3ff: y = 16'h1ed;
			16'h400: y = 16'h1ed;
			16'h401: y = 16'h1ed;
			16'h402: y = 16'h1ed;
			16'h403: y = 16'h1ed;
			16'h404: y = 16'h1ed;
			16'h405: y = 16'h1ed;
			16'h406: y = 16'h1ee;
			16'h407: y = 16'h1ee;
			16'h408: y = 16'h1ee;
			16'h409: y = 16'h1ee;
			16'h40a: y = 16'h1ee;
			16'h40b: y = 16'h1ee;
			16'h40c: y = 16'h1ee;
			16'h40d: y = 16'h1ee;
			16'h40e: y = 16'h1ee;
			16'h40f: y = 16'h1ee;
			16'h410: y = 16'h1ee;
			16'h411: y = 16'h1ee;
			16'h412: y = 16'h1ee;
			16'h413: y = 16'h1ee;
			16'h414: y = 16'h1ee;
			16'h415: y = 16'h1ef;
			16'h416: y = 16'h1ef;
			16'h417: y = 16'h1ef;
			16'h418: y = 16'h1ef;
			16'h419: y = 16'h1ef;
			16'h41a: y = 16'h1ef;
			16'h41b: y = 16'h1ef;
			16'h41c: y = 16'h1ef;
			16'h41d: y = 16'h1ef;
			16'h41e: y = 16'h1ef;
			16'h41f: y = 16'h1ef;
			16'h420: y = 16'h1ef;
			16'h421: y = 16'h1ef;
			16'h422: y = 16'h1ef;
			16'h423: y = 16'h1ef;
			16'h424: y = 16'h1ef;
			16'h425: y = 16'h1f0;
			16'h426: y = 16'h1f0;
			16'h427: y = 16'h1f0;
			16'h428: y = 16'h1f0;
			16'h429: y = 16'h1f0;
			16'h42a: y = 16'h1f0;
			16'h42b: y = 16'h1f0;
			16'h42c: y = 16'h1f0;
			16'h42d: y = 16'h1f0;
			16'h42e: y = 16'h1f0;
			16'h42f: y = 16'h1f0;
			16'h430: y = 16'h1f0;
			16'h431: y = 16'h1f0;
			16'h432: y = 16'h1f0;
			16'h433: y = 16'h1f0;
			16'h434: y = 16'h1f0;
			16'h435: y = 16'h1f0;
			16'h436: y = 16'h1f1;
			16'h437: y = 16'h1f1;
			16'h438: y = 16'h1f1;
			16'h439: y = 16'h1f1;
			16'h43a: y = 16'h1f1;
			16'h43b: y = 16'h1f1;
			16'h43c: y = 16'h1f1;
			16'h43d: y = 16'h1f1;
			16'h43e: y = 16'h1f1;
			16'h43f: y = 16'h1f1;
			16'h440: y = 16'h1f1;
			16'h441: y = 16'h1f1;
			16'h442: y = 16'h1f1;
			16'h443: y = 16'h1f1;
			16'h444: y = 16'h1f1;
			16'h445: y = 16'h1f1;
			16'h446: y = 16'h1f1;
			16'h447: y = 16'h1f1;
			16'h448: y = 16'h1f2;
			16'h449: y = 16'h1f2;
			16'h44a: y = 16'h1f2;
			16'h44b: y = 16'h1f2;
			16'h44c: y = 16'h1f2;
			16'h44d: y = 16'h1f2;
			16'h44e: y = 16'h1f2;
			16'h44f: y = 16'h1f2;
			16'h450: y = 16'h1f2;
			16'h451: y = 16'h1f2;
			16'h452: y = 16'h1f2;
			16'h453: y = 16'h1f2;
			16'h454: y = 16'h1f2;
			16'h455: y = 16'h1f2;
			16'h456: y = 16'h1f2;
			16'h457: y = 16'h1f2;
			16'h458: y = 16'h1f2;
			16'h459: y = 16'h1f2;
			16'h45a: y = 16'h1f2;
			16'h45b: y = 16'h1f3;
			16'h45c: y = 16'h1f3;
			16'h45d: y = 16'h1f3;
			16'h45e: y = 16'h1f3;
			16'h45f: y = 16'h1f3;
			16'h460: y = 16'h1f3;
			16'h461: y = 16'h1f3;
			16'h462: y = 16'h1f3;
			16'h463: y = 16'h1f3;
			16'h464: y = 16'h1f3;
			16'h465: y = 16'h1f3;
			16'h466: y = 16'h1f3;
			16'h467: y = 16'h1f3;
			16'h468: y = 16'h1f3;
			16'h469: y = 16'h1f3;
			16'h46a: y = 16'h1f3;
			16'h46b: y = 16'h1f3;
			16'h46c: y = 16'h1f3;
			16'h46d: y = 16'h1f3;
			16'h46e: y = 16'h1f3;
			16'h46f: y = 16'h1f3;
			16'h470: y = 16'h1f4;
			16'h471: y = 16'h1f4;
			16'h472: y = 16'h1f4;
			16'h473: y = 16'h1f4;
			16'h474: y = 16'h1f4;
			16'h475: y = 16'h1f4;
			16'h476: y = 16'h1f4;
			16'h477: y = 16'h1f4;
			16'h478: y = 16'h1f4;
			16'h479: y = 16'h1f4;
			16'h47a: y = 16'h1f4;
			16'h47b: y = 16'h1f4;
			16'h47c: y = 16'h1f4;
			16'h47d: y = 16'h1f4;
			16'h47e: y = 16'h1f4;
			16'h47f: y = 16'h1f4;
			16'h480: y = 16'h1f4;
			16'h481: y = 16'h1f4;
			16'h482: y = 16'h1f4;
			16'h483: y = 16'h1f4;
			16'h484: y = 16'h1f4;
			16'h485: y = 16'h1f4;
			16'h486: y = 16'h1f5;
			16'h487: y = 16'h1f5;
			16'h488: y = 16'h1f5;
			16'h489: y = 16'h1f5;
			16'h48a: y = 16'h1f5;
			16'h48b: y = 16'h1f5;
			16'h48c: y = 16'h1f5;
			16'h48d: y = 16'h1f5;
			16'h48e: y = 16'h1f5;
			16'h48f: y = 16'h1f5;
			16'h490: y = 16'h1f5;
			16'h491: y = 16'h1f5;
			16'h492: y = 16'h1f5;
			16'h493: y = 16'h1f5;
			16'h494: y = 16'h1f5;
			16'h495: y = 16'h1f5;
			16'h496: y = 16'h1f5;
			16'h497: y = 16'h1f5;
			16'h498: y = 16'h1f5;
			16'h499: y = 16'h1f5;
			16'h49a: y = 16'h1f5;
			16'h49b: y = 16'h1f5;
			16'h49c: y = 16'h1f5;
			16'h49d: y = 16'h1f5;
			16'h49e: y = 16'h1f5;
			16'h49f: y = 16'h1f6;
			16'h4a0: y = 16'h1f6;
			16'h4a1: y = 16'h1f6;
			16'h4a2: y = 16'h1f6;
			16'h4a3: y = 16'h1f6;
			16'h4a4: y = 16'h1f6;
			16'h4a5: y = 16'h1f6;
			16'h4a6: y = 16'h1f6;
			16'h4a7: y = 16'h1f6;
			16'h4a8: y = 16'h1f6;
			16'h4a9: y = 16'h1f6;
			16'h4aa: y = 16'h1f6;
			16'h4ab: y = 16'h1f6;
			16'h4ac: y = 16'h1f6;
			16'h4ad: y = 16'h1f6;
			16'h4ae: y = 16'h1f6;
			16'h4af: y = 16'h1f6;
			16'h4b0: y = 16'h1f6;
			16'h4b1: y = 16'h1f6;
			16'h4b2: y = 16'h1f6;
			16'h4b3: y = 16'h1f6;
			16'h4b4: y = 16'h1f6;
			16'h4b5: y = 16'h1f6;
			16'h4b6: y = 16'h1f6;
			16'h4b7: y = 16'h1f6;
			16'h4b8: y = 16'h1f6;
			16'h4b9: y = 16'h1f6;
			16'h4ba: y = 16'h1f7;
			16'h4bb: y = 16'h1f7;
			16'h4bc: y = 16'h1f7;
			16'h4bd: y = 16'h1f7;
			16'h4be: y = 16'h1f7;
			16'h4bf: y = 16'h1f7;
			16'h4c0: y = 16'h1f7;
			16'h4c1: y = 16'h1f7;
			16'h4c2: y = 16'h1f7;
			16'h4c3: y = 16'h1f7;
			16'h4c4: y = 16'h1f7;
			16'h4c5: y = 16'h1f7;
			16'h4c6: y = 16'h1f7;
			16'h4c7: y = 16'h1f7;
			16'h4c8: y = 16'h1f7;
			16'h4c9: y = 16'h1f7;
			16'h4ca: y = 16'h1f7;
			16'h4cb: y = 16'h1f7;
			16'h4cc: y = 16'h1f7;
			16'h4cd: y = 16'h1f7;
			16'h4ce: y = 16'h1f7;
			16'h4cf: y = 16'h1f7;
			16'h4d0: y = 16'h1f7;
			16'h4d1: y = 16'h1f7;
			16'h4d2: y = 16'h1f7;
			16'h4d3: y = 16'h1f7;
			16'h4d4: y = 16'h1f7;
			16'h4d5: y = 16'h1f7;
			16'h4d6: y = 16'h1f7;
			16'h4d7: y = 16'h1f7;
			16'h4d8: y = 16'h1f7;
			16'h4d9: y = 16'h1f8;
			16'h4da: y = 16'h1f8;
			16'h4db: y = 16'h1f8;
			16'h4dc: y = 16'h1f8;
			16'h4dd: y = 16'h1f8;
			16'h4de: y = 16'h1f8;
			16'h4df: y = 16'h1f8;
			16'h4e0: y = 16'h1f8;
			16'h4e1: y = 16'h1f8;
			16'h4e2: y = 16'h1f8;
			16'h4e3: y = 16'h1f8;
			16'h4e4: y = 16'h1f8;
			16'h4e5: y = 16'h1f8;
			16'h4e6: y = 16'h1f8;
			16'h4e7: y = 16'h1f8;
			16'h4e8: y = 16'h1f8;
			16'h4e9: y = 16'h1f8;
			16'h4ea: y = 16'h1f8;
			16'h4eb: y = 16'h1f8;
			16'h4ec: y = 16'h1f8;
			16'h4ed: y = 16'h1f8;
			16'h4ee: y = 16'h1f8;
			16'h4ef: y = 16'h1f8;
			16'h4f0: y = 16'h1f8;
			16'h4f1: y = 16'h1f8;
			16'h4f2: y = 16'h1f8;
			16'h4f3: y = 16'h1f8;
			16'h4f4: y = 16'h1f8;
			16'h4f5: y = 16'h1f8;
			16'h4f6: y = 16'h1f8;
			16'h4f7: y = 16'h1f8;
			16'h4f8: y = 16'h1f8;
			16'h4f9: y = 16'h1f8;
			16'h4fa: y = 16'h1f8;
			16'h4fb: y = 16'h1f9;
			16'h4fc: y = 16'h1f9;
			16'h4fd: y = 16'h1f9;
			16'h4fe: y = 16'h1f9;
			16'h4ff: y = 16'h1f9;
			16'h500: y = 16'h1f9;
			16'h501: y = 16'h1f9;
			16'h502: y = 16'h1f9;
			16'h503: y = 16'h1f9;
			16'h504: y = 16'h1f9;
			16'h505: y = 16'h1f9;
			16'h506: y = 16'h1f9;
			16'h507: y = 16'h1f9;
			16'h508: y = 16'h1f9;
			16'h509: y = 16'h1f9;
			16'h50a: y = 16'h1f9;
			16'h50b: y = 16'h1f9;
			16'h50c: y = 16'h1f9;
			16'h50d: y = 16'h1f9;
			16'h50e: y = 16'h1f9;
			16'h50f: y = 16'h1f9;
			16'h510: y = 16'h1f9;
			16'h511: y = 16'h1f9;
			16'h512: y = 16'h1f9;
			16'h513: y = 16'h1f9;
			16'h514: y = 16'h1f9;
			16'h515: y = 16'h1f9;
			16'h516: y = 16'h1f9;
			16'h517: y = 16'h1f9;
			16'h518: y = 16'h1f9;
			16'h519: y = 16'h1f9;
			16'h51a: y = 16'h1f9;
			16'h51b: y = 16'h1f9;
			16'h51c: y = 16'h1f9;
			16'h51d: y = 16'h1f9;
			16'h51e: y = 16'h1f9;
			16'h51f: y = 16'h1f9;
			16'h520: y = 16'h1f9;
			16'h521: y = 16'h1f9;
			16'h522: y = 16'h1f9;
			16'h523: y = 16'h1fa;
			16'h524: y = 16'h1fa;
			16'h525: y = 16'h1fa;
			16'h526: y = 16'h1fa;
			16'h527: y = 16'h1fa;
			16'h528: y = 16'h1fa;
			16'h529: y = 16'h1fa;
			16'h52a: y = 16'h1fa;
			16'h52b: y = 16'h1fa;
			16'h52c: y = 16'h1fa;
			16'h52d: y = 16'h1fa;
			16'h52e: y = 16'h1fa;
			16'h52f: y = 16'h1fa;
			16'h530: y = 16'h1fa;
			16'h531: y = 16'h1fa;
			16'h532: y = 16'h1fa;
			16'h533: y = 16'h1fa;
			16'h534: y = 16'h1fa;
			16'h535: y = 16'h1fa;
			16'h536: y = 16'h1fa;
			16'h537: y = 16'h1fa;
			16'h538: y = 16'h1fa;
			16'h539: y = 16'h1fa;
			16'h53a: y = 16'h1fa;
			16'h53b: y = 16'h1fa;
			16'h53c: y = 16'h1fa;
			16'h53d: y = 16'h1fa;
			16'h53e: y = 16'h1fa;
			16'h53f: y = 16'h1fa;
			16'h540: y = 16'h1fa;
			16'h541: y = 16'h1fa;
			16'h542: y = 16'h1fa;
			16'h543: y = 16'h1fa;
			16'h544: y = 16'h1fa;
			16'h545: y = 16'h1fa;
			16'h546: y = 16'h1fa;
			16'h547: y = 16'h1fa;
			16'h548: y = 16'h1fa;
			16'h549: y = 16'h1fa;
			16'h54a: y = 16'h1fa;
			16'h54b: y = 16'h1fa;
			16'h54c: y = 16'h1fa;
			16'h54d: y = 16'h1fa;
			16'h54e: y = 16'h1fa;
			16'h54f: y = 16'h1fa;
			16'h550: y = 16'h1fa;
			16'h551: y = 16'h1fa;
			16'h552: y = 16'h1fb;
			16'h553: y = 16'h1fb;
			16'h554: y = 16'h1fb;
			16'h555: y = 16'h1fb;
			16'h556: y = 16'h1fb;
			16'h557: y = 16'h1fb;
			16'h558: y = 16'h1fb;
			16'h559: y = 16'h1fb;
			16'h55a: y = 16'h1fb;
			16'h55b: y = 16'h1fb;
			16'h55c: y = 16'h1fb;
			16'h55d: y = 16'h1fb;
			16'h55e: y = 16'h1fb;
			16'h55f: y = 16'h1fb;
			16'h560: y = 16'h1fb;
			16'h561: y = 16'h1fb;
			16'h562: y = 16'h1fb;
			16'h563: y = 16'h1fb;
			16'h564: y = 16'h1fb;
			16'h565: y = 16'h1fb;
			16'h566: y = 16'h1fb;
			16'h567: y = 16'h1fb;
			16'h568: y = 16'h1fb;
			16'h569: y = 16'h1fb;
			16'h56a: y = 16'h1fb;
			16'h56b: y = 16'h1fb;
			16'h56c: y = 16'h1fb;
			16'h56d: y = 16'h1fb;
			16'h56e: y = 16'h1fb;
			16'h56f: y = 16'h1fb;
			16'h570: y = 16'h1fb;
			16'h571: y = 16'h1fb;
			16'h572: y = 16'h1fb;
			16'h573: y = 16'h1fb;
			16'h574: y = 16'h1fb;
			16'h575: y = 16'h1fb;
			16'h576: y = 16'h1fb;
			16'h577: y = 16'h1fb;
			16'h578: y = 16'h1fb;
			16'h579: y = 16'h1fb;
			16'h57a: y = 16'h1fb;
			16'h57b: y = 16'h1fb;
			16'h57c: y = 16'h1fb;
			16'h57d: y = 16'h1fb;
			16'h57e: y = 16'h1fb;
			16'h57f: y = 16'h1fb;
			16'h580: y = 16'h1fb;
			16'h581: y = 16'h1fb;
			16'h582: y = 16'h1fb;
			16'h583: y = 16'h1fb;
			16'h584: y = 16'h1fb;
			16'h585: y = 16'h1fb;
			16'h586: y = 16'h1fb;
			16'h587: y = 16'h1fb;
			16'h588: y = 16'h1fb;
			16'h589: y = 16'h1fb;
			16'h58a: y = 16'h1fb;
			16'h58b: y = 16'h1fc;
			16'h58c: y = 16'h1fc;
			16'h58d: y = 16'h1fc;
			16'h58e: y = 16'h1fc;
			16'h58f: y = 16'h1fc;
			16'h590: y = 16'h1fc;
			16'h591: y = 16'h1fc;
			16'h592: y = 16'h1fc;
			16'h593: y = 16'h1fc;
			16'h594: y = 16'h1fc;
			16'h595: y = 16'h1fc;
			16'h596: y = 16'h1fc;
			16'h597: y = 16'h1fc;
			16'h598: y = 16'h1fc;
			16'h599: y = 16'h1fc;
			16'h59a: y = 16'h1fc;
			16'h59b: y = 16'h1fc;
			16'h59c: y = 16'h1fc;
			16'h59d: y = 16'h1fc;
			16'h59e: y = 16'h1fc;
			16'h59f: y = 16'h1fc;
			16'h5a0: y = 16'h1fc;
			16'h5a1: y = 16'h1fc;
			16'h5a2: y = 16'h1fc;
			16'h5a3: y = 16'h1fc;
			16'h5a4: y = 16'h1fc;
			16'h5a5: y = 16'h1fc;
			16'h5a6: y = 16'h1fc;
			16'h5a7: y = 16'h1fc;
			16'h5a8: y = 16'h1fc;
			16'h5a9: y = 16'h1fc;
			16'h5aa: y = 16'h1fc;
			16'h5ab: y = 16'h1fc;
			16'h5ac: y = 16'h1fc;
			16'h5ad: y = 16'h1fc;
			16'h5ae: y = 16'h1fc;
			16'h5af: y = 16'h1fc;
			16'h5b0: y = 16'h1fc;
			16'h5b1: y = 16'h1fc;
			16'h5b2: y = 16'h1fc;
			16'h5b3: y = 16'h1fc;
			16'h5b4: y = 16'h1fc;
			16'h5b5: y = 16'h1fc;
			16'h5b6: y = 16'h1fc;
			16'h5b7: y = 16'h1fc;
			16'h5b8: y = 16'h1fc;
			16'h5b9: y = 16'h1fc;
			16'h5ba: y = 16'h1fc;
			16'h5bb: y = 16'h1fc;
			16'h5bc: y = 16'h1fc;
			16'h5bd: y = 16'h1fc;
			16'h5be: y = 16'h1fc;
			16'h5bf: y = 16'h1fc;
			16'h5c0: y = 16'h1fc;
			16'h5c1: y = 16'h1fc;
			16'h5c2: y = 16'h1fc;
			16'h5c3: y = 16'h1fc;
			16'h5c4: y = 16'h1fc;
			16'h5c5: y = 16'h1fc;
			16'h5c6: y = 16'h1fc;
			16'h5c7: y = 16'h1fc;
			16'h5c8: y = 16'h1fc;
			16'h5c9: y = 16'h1fc;
			16'h5ca: y = 16'h1fc;
			16'h5cb: y = 16'h1fc;
			16'h5cc: y = 16'h1fc;
			16'h5cd: y = 16'h1fc;
			16'h5ce: y = 16'h1fc;
			16'h5cf: y = 16'h1fc;
			16'h5d0: y = 16'h1fc;
			16'h5d1: y = 16'h1fc;
			16'h5d2: y = 16'h1fc;
			16'h5d3: y = 16'h1fc;
			16'h5d4: y = 16'h1fc;
			16'h5d5: y = 16'h1fd;
			16'h5d6: y = 16'h1fd;
			16'h5d7: y = 16'h1fd;
			16'h5d8: y = 16'h1fd;
			16'h5d9: y = 16'h1fd;
			16'h5da: y = 16'h1fd;
			16'h5db: y = 16'h1fd;
			16'h5dc: y = 16'h1fd;
			16'h5dd: y = 16'h1fd;
			16'h5de: y = 16'h1fd;
			16'h5df: y = 16'h1fd;
			16'h5e0: y = 16'h1fd;
			16'h5e1: y = 16'h1fd;
			16'h5e2: y = 16'h1fd;
			16'h5e3: y = 16'h1fd;
			16'h5e4: y = 16'h1fd;
			16'h5e5: y = 16'h1fd;
			16'h5e6: y = 16'h1fd;
			16'h5e7: y = 16'h1fd;
			16'h5e8: y = 16'h1fd;
			16'h5e9: y = 16'h1fd;
			16'h5ea: y = 16'h1fd;
			16'h5eb: y = 16'h1fd;
			16'h5ec: y = 16'h1fd;
			16'h5ed: y = 16'h1fd;
			16'h5ee: y = 16'h1fd;
			16'h5ef: y = 16'h1fd;
			16'h5f0: y = 16'h1fd;
			16'h5f1: y = 16'h1fd;
			16'h5f2: y = 16'h1fd;
			16'h5f3: y = 16'h1fd;
			16'h5f4: y = 16'h1fd;
			16'h5f5: y = 16'h1fd;
			16'h5f6: y = 16'h1fd;
			16'h5f7: y = 16'h1fd;
			16'h5f8: y = 16'h1fd;
			16'h5f9: y = 16'h1fd;
			16'h5fa: y = 16'h1fd;
			16'h5fb: y = 16'h1fd;
			16'h5fc: y = 16'h1fd;
			16'h5fd: y = 16'h1fd;
			16'h5fe: y = 16'h1fd;
			16'h5ff: y = 16'h1fd;
			16'h600: y = 16'h1fd;
			16'h601: y = 16'h1fd;
			16'h602: y = 16'h1fd;
			16'h603: y = 16'h1fd;
			16'h604: y = 16'h1fd;
			16'h605: y = 16'h1fd;
			16'h606: y = 16'h1fd;
			16'h607: y = 16'h1fd;
			16'h608: y = 16'h1fd;
			16'h609: y = 16'h1fd;
			16'h60a: y = 16'h1fd;
			16'h60b: y = 16'h1fd;
			16'h60c: y = 16'h1fd;
			16'h60d: y = 16'h1fd;
			16'h60e: y = 16'h1fd;
			16'h60f: y = 16'h1fd;
			16'h610: y = 16'h1fd;
			16'h611: y = 16'h1fd;
			16'h612: y = 16'h1fd;
			16'h613: y = 16'h1fd;
			16'h614: y = 16'h1fd;
			16'h615: y = 16'h1fd;
			16'h616: y = 16'h1fd;
			16'h617: y = 16'h1fd;
			16'h618: y = 16'h1fd;
			16'h619: y = 16'h1fd;
			16'h61a: y = 16'h1fd;
			16'h61b: y = 16'h1fd;
			16'h61c: y = 16'h1fd;
			16'h61d: y = 16'h1fd;
			16'h61e: y = 16'h1fd;
			16'h61f: y = 16'h1fd;
			16'h620: y = 16'h1fd;
			16'h621: y = 16'h1fd;
			16'h622: y = 16'h1fd;
			16'h623: y = 16'h1fd;
			16'h624: y = 16'h1fd;
			16'h625: y = 16'h1fd;
			16'h626: y = 16'h1fd;
			16'h627: y = 16'h1fd;
			16'h628: y = 16'h1fd;
			16'h629: y = 16'h1fd;
			16'h62a: y = 16'h1fd;
			16'h62b: y = 16'h1fd;
			16'h62c: y = 16'h1fd;
			16'h62d: y = 16'h1fd;
			16'h62e: y = 16'h1fd;
			16'h62f: y = 16'h1fd;
			16'h630: y = 16'h1fd;
			16'h631: y = 16'h1fd;
			16'h632: y = 16'h1fd;
			16'h633: y = 16'h1fd;
			16'h634: y = 16'h1fd;
			16'h635: y = 16'h1fd;
			16'h636: y = 16'h1fd;
			16'h637: y = 16'h1fd;
			16'h638: y = 16'h1fd;
			16'h639: y = 16'h1fd;
			16'h63a: y = 16'h1fd;
			16'h63b: y = 16'h1fd;
			16'h63c: y = 16'h1fd;
			16'h63d: y = 16'h1fe;
			16'h63e: y = 16'h1fe;
			16'h63f: y = 16'h1fe;
			16'h640: y = 16'h1fe;
			16'h641: y = 16'h1fe;
			16'h642: y = 16'h1fe;
			16'h643: y = 16'h1fe;
			16'h644: y = 16'h1fe;
			16'h645: y = 16'h1fe;
			16'h646: y = 16'h1fe;
			16'h647: y = 16'h1fe;
			16'h648: y = 16'h1fe;
			16'h649: y = 16'h1fe;
			16'h64a: y = 16'h1fe;
			16'h64b: y = 16'h1fe;
			16'h64c: y = 16'h1fe;
			16'h64d: y = 16'h1fe;
			16'h64e: y = 16'h1fe;
			16'h64f: y = 16'h1fe;
			16'h650: y = 16'h1fe;
			16'h651: y = 16'h1fe;
			16'h652: y = 16'h1fe;
			16'h653: y = 16'h1fe;
			16'h654: y = 16'h1fe;
			16'h655: y = 16'h1fe;
			16'h656: y = 16'h1fe;
			16'h657: y = 16'h1fe;
			16'h658: y = 16'h1fe;
			16'h659: y = 16'h1fe;
			16'h65a: y = 16'h1fe;
			16'h65b: y = 16'h1fe;
			16'h65c: y = 16'h1fe;
			16'h65d: y = 16'h1fe;
			16'h65e: y = 16'h1fe;
			16'h65f: y = 16'h1fe;
			16'h660: y = 16'h1fe;
			16'h661: y = 16'h1fe;
			16'h662: y = 16'h1fe;
			16'h663: y = 16'h1fe;
			16'h664: y = 16'h1fe;
			16'h665: y = 16'h1fe;
			16'h666: y = 16'h1fe;
			16'h667: y = 16'h1fe;
			16'h668: y = 16'h1fe;
			16'h669: y = 16'h1fe;
			16'h66a: y = 16'h1fe;
			16'h66b: y = 16'h1fe;
			16'h66c: y = 16'h1fe;
			16'h66d: y = 16'h1fe;
			16'h66e: y = 16'h1fe;
			16'h66f: y = 16'h1fe;
			16'h670: y = 16'h1fe;
			16'h671: y = 16'h1fe;
			16'h672: y = 16'h1fe;
			16'h673: y = 16'h1fe;
			16'h674: y = 16'h1fe;
			16'h675: y = 16'h1fe;
			16'h676: y = 16'h1fe;
			16'h677: y = 16'h1fe;
			16'h678: y = 16'h1fe;
			16'h679: y = 16'h1fe;
			16'h67a: y = 16'h1fe;
			16'h67b: y = 16'h1fe;
			16'h67c: y = 16'h1fe;
			16'h67d: y = 16'h1fe;
			16'h67e: y = 16'h1fe;
			16'h67f: y = 16'h1fe;
			16'h680: y = 16'h1fe;
			16'h681: y = 16'h1fe;
			16'h682: y = 16'h1fe;
			16'h683: y = 16'h1fe;
			16'h684: y = 16'h1fe;
			16'h685: y = 16'h1fe;
			16'h686: y = 16'h1fe;
			16'h687: y = 16'h1fe;
			16'h688: y = 16'h1fe;
			16'h689: y = 16'h1fe;
			16'h68a: y = 16'h1fe;
			16'h68b: y = 16'h1fe;
			16'h68c: y = 16'h1fe;
			16'h68d: y = 16'h1fe;
			16'h68e: y = 16'h1fe;
			16'h68f: y = 16'h1fe;
			16'h690: y = 16'h1fe;
			16'h691: y = 16'h1fe;
			16'h692: y = 16'h1fe;
			16'h693: y = 16'h1fe;
			16'h694: y = 16'h1fe;
			16'h695: y = 16'h1fe;
			16'h696: y = 16'h1fe;
			16'h697: y = 16'h1fe;
			16'h698: y = 16'h1fe;
			16'h699: y = 16'h1fe;
			16'h69a: y = 16'h1fe;
			16'h69b: y = 16'h1fe;
			16'h69c: y = 16'h1fe;
			16'h69d: y = 16'h1fe;
			16'h69e: y = 16'h1fe;
			16'h69f: y = 16'h1fe;
			16'h6a0: y = 16'h1fe;
			16'h6a1: y = 16'h1fe;
			16'h6a2: y = 16'h1fe;
			16'h6a3: y = 16'h1fe;
			16'h6a4: y = 16'h1fe;
			16'h6a5: y = 16'h1fe;
			16'h6a6: y = 16'h1fe;
			16'h6a7: y = 16'h1fe;
			16'h6a8: y = 16'h1fe;
			16'h6a9: y = 16'h1fe;
			16'h6aa: y = 16'h1fe;
			16'h6ab: y = 16'h1fe;
			16'h6ac: y = 16'h1fe;
			16'h6ad: y = 16'h1fe;
			16'h6ae: y = 16'h1fe;
			16'h6af: y = 16'h1fe;
			16'h6b0: y = 16'h1fe;
			16'h6b1: y = 16'h1fe;
			16'h6b2: y = 16'h1fe;
			16'h6b3: y = 16'h1fe;
			16'h6b4: y = 16'h1fe;
			16'h6b5: y = 16'h1fe;
			16'h6b6: y = 16'h1fe;
			16'h6b7: y = 16'h1fe;
			16'h6b8: y = 16'h1fe;
			16'h6b9: y = 16'h1fe;
			16'h6ba: y = 16'h1fe;
			16'h6bb: y = 16'h1fe;
			16'h6bc: y = 16'h1fe;
			16'h6bd: y = 16'h1fe;
			16'h6be: y = 16'h1fe;
			16'h6bf: y = 16'h1fe;
			16'h6c0: y = 16'h1fe;
			16'h6c1: y = 16'h1fe;
			16'h6c2: y = 16'h1fe;
			16'h6c3: y = 16'h1fe;
			16'h6c4: y = 16'h1fe;
			16'h6c5: y = 16'h1fe;
			16'h6c6: y = 16'h1fe;
			16'h6c7: y = 16'h1fe;
			16'h6c8: y = 16'h1fe;
			16'h6c9: y = 16'h1fe;
			16'h6ca: y = 16'h1fe;
			16'h6cb: y = 16'h1fe;
			16'h6cc: y = 16'h1fe;
			16'h6cd: y = 16'h1fe;
			16'h6ce: y = 16'h1fe;
			16'h6cf: y = 16'h1fe;
			16'h6d0: y = 16'h1fe;
			16'h6d1: y = 16'h1fe;
			16'h6d2: y = 16'h1fe;
			16'h6d3: y = 16'h1fe;
			16'h6d4: y = 16'h1fe;
			16'h6d5: y = 16'h1fe;
			16'h6d6: y = 16'h1fe;
			16'h6d7: y = 16'h1fe;
			16'h6d8: y = 16'h1fe;
			16'h6d9: y = 16'h1fe;
			16'h6da: y = 16'h1fe;
			16'h6db: y = 16'h1fe;
			16'h6dc: y = 16'h1fe;
			16'h6dd: y = 16'h1fe;
			16'h6de: y = 16'h1fe;
			16'h6df: y = 16'h1fe;
			16'h6e0: y = 16'h1fe;
			16'h6e1: y = 16'h1fe;
			16'h6e2: y = 16'h1fe;
			16'h6e3: y = 16'h1fe;
			16'h6e4: y = 16'h1fe;
			16'h6e5: y = 16'h1fe;
			16'h6e6: y = 16'h1fe;
			16'h6e7: y = 16'h1fe;
			16'h6e8: y = 16'h1fe;
			16'h6e9: y = 16'h1fe;
			16'h6ea: y = 16'h1fe;
			16'h6eb: y = 16'h1fe;
			16'h6ec: y = 16'h1fe;
			16'h6ed: y = 16'h1fe;
			16'h6ee: y = 16'h1fe;
			16'h6ef: y = 16'h1ff;
			16'h6f0: y = 16'h1ff;
			16'h6f1: y = 16'h1ff;
			16'h6f2: y = 16'h1ff;
			16'h6f3: y = 16'h1ff;
			16'h6f4: y = 16'h1ff;
			16'h6f5: y = 16'h1ff;
			16'h6f6: y = 16'h1ff;
			16'h6f7: y = 16'h1ff;
			16'h6f8: y = 16'h1ff;
			16'h6f9: y = 16'h1ff;
			16'h6fa: y = 16'h1ff;
			16'h6fb: y = 16'h1ff;
			16'h6fc: y = 16'h1ff;
			16'h6fd: y = 16'h1ff;
			16'h6fe: y = 16'h1ff;
			16'h6ff: y = 16'h1ff;
			16'h700: y = 16'h1ff;
			16'h701: y = 16'h1ff;
			16'h702: y = 16'h1ff;
			16'h703: y = 16'h1ff;
			16'h704: y = 16'h1ff;
			16'h705: y = 16'h1ff;
			16'h706: y = 16'h1ff;
			16'h707: y = 16'h1ff;
			16'h708: y = 16'h1ff;
			16'h709: y = 16'h1ff;
			16'h70a: y = 16'h1ff;
			16'h70b: y = 16'h1ff;
			16'h70c: y = 16'h1ff;
			16'h70d: y = 16'h1ff;
			16'h70e: y = 16'h1ff;
			16'h70f: y = 16'h1ff;
			16'h710: y = 16'h1ff;
			16'h711: y = 16'h1ff;
			16'h712: y = 16'h1ff;
			16'h713: y = 16'h1ff;
			16'h714: y = 16'h1ff;
			16'h715: y = 16'h1ff;
			16'h716: y = 16'h1ff;
			16'h717: y = 16'h1ff;
			16'h718: y = 16'h1ff;
			16'h719: y = 16'h1ff;
			16'h71a: y = 16'h1ff;
			16'h71b: y = 16'h1ff;
			16'h71c: y = 16'h1ff;
			16'h71d: y = 16'h1ff;
			16'h71e: y = 16'h1ff;
			16'h71f: y = 16'h1ff;
			16'h720: y = 16'h1ff;
			16'h721: y = 16'h1ff;
			16'h722: y = 16'h1ff;
			16'h723: y = 16'h1ff;
			16'h724: y = 16'h1ff;
			16'h725: y = 16'h1ff;
			16'h726: y = 16'h1ff;
			16'h727: y = 16'h1ff;
			16'h728: y = 16'h1ff;
			16'h729: y = 16'h1ff;
			16'h72a: y = 16'h1ff;
			16'h72b: y = 16'h1ff;
			16'h72c: y = 16'h1ff;
			16'h72d: y = 16'h1ff;
			16'h72e: y = 16'h1ff;
			16'h72f: y = 16'h1ff;
			16'h730: y = 16'h1ff;
			16'h731: y = 16'h1ff;
			16'h732: y = 16'h1ff;
			16'h733: y = 16'h1ff;
			16'h734: y = 16'h1ff;
			16'h735: y = 16'h1ff;
			16'h736: y = 16'h1ff;
			16'h737: y = 16'h1ff;
			16'h738: y = 16'h1ff;
			16'h739: y = 16'h1ff;
			16'h73a: y = 16'h1ff;
			16'h73b: y = 16'h1ff;
			16'h73c: y = 16'h1ff;
			16'h73d: y = 16'h1ff;
			16'h73e: y = 16'h1ff;
			16'h73f: y = 16'h1ff;
			16'h740: y = 16'h1ff;
			16'h741: y = 16'h1ff;
			16'h742: y = 16'h1ff;
			16'h743: y = 16'h1ff;
			16'h744: y = 16'h1ff;
			16'h745: y = 16'h1ff;
			16'h746: y = 16'h1ff;
			16'h747: y = 16'h1ff;
			16'h748: y = 16'h1ff;
			16'h749: y = 16'h1ff;
			16'h74a: y = 16'h1ff;
			16'h74b: y = 16'h1ff;
			16'h74c: y = 16'h1ff;
			16'h74d: y = 16'h1ff;
			16'h74e: y = 16'h1ff;
			16'h74f: y = 16'h1ff;
			16'h750: y = 16'h1ff;
			16'h751: y = 16'h1ff;
			16'h752: y = 16'h1ff;
			16'h753: y = 16'h1ff;
			16'h754: y = 16'h1ff;
			16'h755: y = 16'h1ff;
			16'h756: y = 16'h1ff;
			16'h757: y = 16'h1ff;
			16'h758: y = 16'h1ff;
			16'h759: y = 16'h1ff;
			16'h75a: y = 16'h1ff;
			16'h75b: y = 16'h1ff;
			16'h75c: y = 16'h1ff;
			16'h75d: y = 16'h1ff;
			16'h75e: y = 16'h1ff;
			16'h75f: y = 16'h1ff;
			16'h760: y = 16'h1ff;
			16'h761: y = 16'h1ff;
			16'h762: y = 16'h1ff;
			16'h763: y = 16'h1ff;
			16'h764: y = 16'h1ff;
			16'h765: y = 16'h1ff;
			16'h766: y = 16'h1ff;
			16'h767: y = 16'h1ff;
			16'h768: y = 16'h1ff;
			16'h769: y = 16'h1ff;
			16'h76a: y = 16'h1ff;
			16'h76b: y = 16'h1ff;
			16'h76c: y = 16'h1ff;
			16'h76d: y = 16'h1ff;
			16'h76e: y = 16'h1ff;
			16'h76f: y = 16'h1ff;
			16'h770: y = 16'h1ff;
			16'h771: y = 16'h1ff;
			16'h772: y = 16'h1ff;
			16'h773: y = 16'h1ff;
			16'h774: y = 16'h1ff;
			16'h775: y = 16'h1ff;
			16'h776: y = 16'h1ff;
			16'h777: y = 16'h1ff;
			16'h778: y = 16'h1ff;
			16'h779: y = 16'h1ff;
			16'h77a: y = 16'h1ff;
			16'h77b: y = 16'h1ff;
			16'h77c: y = 16'h1ff;
			16'h77d: y = 16'h1ff;
			16'h77e: y = 16'h1ff;
			16'h77f: y = 16'h1ff;
			16'h780: y = 16'h1ff;
			16'h781: y = 16'h1ff;
			16'h782: y = 16'h1ff;
			16'h783: y = 16'h1ff;
			16'h784: y = 16'h1ff;
			16'h785: y = 16'h1ff;
			16'h786: y = 16'h1ff;
			16'h787: y = 16'h1ff;
			16'h788: y = 16'h1ff;
			16'h789: y = 16'h1ff;
			16'h78a: y = 16'h1ff;
			16'h78b: y = 16'h1ff;
			16'h78c: y = 16'h1ff;
			16'h78d: y = 16'h1ff;
			16'h78e: y = 16'h1ff;
			16'h78f: y = 16'h1ff;
			16'h790: y = 16'h1ff;
			16'h791: y = 16'h1ff;
			16'h792: y = 16'h1ff;
			16'h793: y = 16'h1ff;
			16'h794: y = 16'h1ff;
			16'h795: y = 16'h1ff;
			16'h796: y = 16'h1ff;
			16'h797: y = 16'h1ff;
			16'h798: y = 16'h1ff;
			16'h799: y = 16'h1ff;
			16'h79a: y = 16'h1ff;
			16'h79b: y = 16'h1ff;
			16'h79c: y = 16'h1ff;
			16'h79d: y = 16'h1ff;
			16'h79e: y = 16'h1ff;
			16'h79f: y = 16'h1ff;
			16'h7a0: y = 16'h1ff;
			16'h7a1: y = 16'h1ff;
			16'h7a2: y = 16'h1ff;
			16'h7a3: y = 16'h1ff;
			16'h7a4: y = 16'h1ff;
			16'h7a5: y = 16'h1ff;
			16'h7a6: y = 16'h1ff;
			16'h7a7: y = 16'h1ff;
			16'h7a8: y = 16'h1ff;
			16'h7a9: y = 16'h1ff;
			16'h7aa: y = 16'h1ff;
			16'h7ab: y = 16'h1ff;
			16'h7ac: y = 16'h1ff;
			16'h7ad: y = 16'h1ff;
			16'h7ae: y = 16'h1ff;
			16'h7af: y = 16'h1ff;
			16'h7b0: y = 16'h1ff;
			16'h7b1: y = 16'h1ff;
			16'h7b2: y = 16'h1ff;
			16'h7b3: y = 16'h1ff;
			16'h7b4: y = 16'h1ff;
			16'h7b5: y = 16'h1ff;
			16'h7b6: y = 16'h1ff;
			16'h7b7: y = 16'h1ff;
			16'h7b8: y = 16'h1ff;
			16'h7b9: y = 16'h1ff;
			16'h7ba: y = 16'h1ff;
			16'h7bb: y = 16'h1ff;
			16'h7bc: y = 16'h1ff;
			16'h7bd: y = 16'h1ff;
			16'h7be: y = 16'h1ff;
			16'h7bf: y = 16'h1ff;
			16'h7c0: y = 16'h1ff;
			16'h7c1: y = 16'h1ff;
			16'h7c2: y = 16'h1ff;
			16'h7c3: y = 16'h1ff;
			16'h7c4: y = 16'h1ff;
			16'h7c5: y = 16'h1ff;
			16'h7c6: y = 16'h1ff;
			16'h7c7: y = 16'h1ff;
			16'h7c8: y = 16'h1ff;
			16'h7c9: y = 16'h1ff;
			16'h7ca: y = 16'h1ff;
			16'h7cb: y = 16'h1ff;
			16'h7cc: y = 16'h1ff;
			16'h7cd: y = 16'h1ff;
			16'h7ce: y = 16'h1ff;
			16'h7cf: y = 16'h1ff;
			16'h7d0: y = 16'h1ff;
			16'h7d1: y = 16'h1ff;
			16'h7d2: y = 16'h1ff;
			16'h7d3: y = 16'h1ff;
			16'h7d4: y = 16'h1ff;
			16'h7d5: y = 16'h1ff;
			16'h7d6: y = 16'h1ff;
			16'h7d7: y = 16'h1ff;
			16'h7d8: y = 16'h1ff;
			16'h7d9: y = 16'h1ff;
			16'h7da: y = 16'h1ff;
			16'h7db: y = 16'h1ff;
			16'h7dc: y = 16'h1ff;
			16'h7dd: y = 16'h1ff;
			16'h7de: y = 16'h1ff;
			16'h7df: y = 16'h1ff;
			16'h7e0: y = 16'h1ff;
			16'h7e1: y = 16'h1ff;
			16'h7e2: y = 16'h1ff;
			16'h7e3: y = 16'h1ff;
			16'h7e4: y = 16'h1ff;
			16'h7e5: y = 16'h1ff;
			16'h7e6: y = 16'h1ff;
			16'h7e7: y = 16'h1ff;
			16'h7e8: y = 16'h1ff;
			16'h7e9: y = 16'h1ff;
			16'h7ea: y = 16'h1ff;
			16'h7eb: y = 16'h1ff;
			16'h7ec: y = 16'h1ff;
			16'h7ed: y = 16'h1ff;
			16'h7ee: y = 16'h1ff;
			16'h7ef: y = 16'h1ff;
			16'h7f0: y = 16'h1ff;
			16'h7f1: y = 16'h1ff;
			16'h7f2: y = 16'h1ff;
			16'h7f3: y = 16'h1ff;
			16'h7f4: y = 16'h1ff;
			16'h7f5: y = 16'h1ff;
			16'h7f6: y = 16'h1ff;
			16'h7f7: y = 16'h1ff;
			16'h7f8: y = 16'h1ff;
			16'h7f9: y = 16'h1ff;
			16'h7fa: y = 16'h1ff;
			16'h7fb: y = 16'h1ff;
			16'h7fc: y = 16'h1ff;
			16'h7fd: y = 16'h1ff;
			16'h7fe: y = 16'h1ff;
			16'h7ff: y = 16'h1ff;
			16'h800: y = 16'h1ff;
			16'h801: y = 16'h1ff;
			16'h802: y = 16'h1ff;
			16'h803: y = 16'h1ff;
			16'h804: y = 16'h1ff;
			16'h805: y = 16'h1ff;
			16'h806: y = 16'h1ff;
			16'h807: y = 16'h1ff;
			16'h808: y = 16'h1ff;
			16'h809: y = 16'h1ff;
			16'h80a: y = 16'h1ff;
			16'h80b: y = 16'h1ff;
			16'h80c: y = 16'h1ff;
			16'h80d: y = 16'h1ff;
			16'h80e: y = 16'h1ff;
			16'h80f: y = 16'h1ff;
			16'h810: y = 16'h1ff;
			16'h811: y = 16'h1ff;
			16'h812: y = 16'h1ff;
			16'h813: y = 16'h1ff;
			16'h814: y = 16'h1ff;
			16'h815: y = 16'h1ff;
			16'h816: y = 16'h1ff;
			16'h817: y = 16'h1ff;
			16'h818: y = 16'h1ff;
			16'h819: y = 16'h1ff;
			16'h81a: y = 16'h1ff;
			16'h81b: y = 16'h1ff;
			16'h81c: y = 16'h1ff;
			16'h81d: y = 16'h1ff;
			16'h81e: y = 16'h1ff;
			16'h81f: y = 16'h1ff;
			16'h820: y = 16'h1ff;
			16'h821: y = 16'h1ff;
			16'h822: y = 16'h1ff;
			16'h823: y = 16'h1ff;
			16'h824: y = 16'h1ff;
			16'h825: y = 16'h1ff;
			16'h826: y = 16'h1ff;
			16'h827: y = 16'h1ff;
			16'h828: y = 16'h1ff;
			16'h829: y = 16'h1ff;
			16'h82a: y = 16'h1ff;
			16'h82b: y = 16'h1ff;
			16'h82c: y = 16'h1ff;
			16'h82d: y = 16'h1ff;
			16'h82e: y = 16'h1ff;
			16'h82f: y = 16'h1ff;
			16'h830: y = 16'h1ff;
			16'h831: y = 16'h1ff;
			16'h832: y = 16'h1ff;
			16'h833: y = 16'h1ff;
			16'h834: y = 16'h1ff;
			16'h835: y = 16'h1ff;
			16'h836: y = 16'h1ff;
			16'h837: y = 16'h1ff;
			16'h838: y = 16'h1ff;
			16'h839: y = 16'h1ff;
			16'h83a: y = 16'h1ff;
			16'h83b: y = 16'h1ff;
			16'h83c: y = 16'h1ff;
			16'h83d: y = 16'h1ff;
			16'h83e: y = 16'h1ff;
			16'h83f: y = 16'h1ff;
			16'h840: y = 16'h1ff;
			16'h841: y = 16'h1ff;
			16'h842: y = 16'h1ff;
			16'h843: y = 16'h1ff;
			16'h844: y = 16'h1ff;
			16'h845: y = 16'h1ff;
			16'h846: y = 16'h1ff;
			16'h847: y = 16'h1ff;
			16'h848: y = 16'h1ff;
			16'h849: y = 16'h1ff;
			16'h84a: y = 16'h1ff;
			16'h84b: y = 16'h1ff;
			16'h84c: y = 16'h1ff;
			16'h84d: y = 16'h1ff;
			16'h84e: y = 16'h1ff;
			16'h84f: y = 16'h1ff;
			16'h850: y = 16'h1ff;
			16'h851: y = 16'h1ff;
			16'h852: y = 16'h1ff;
			16'h853: y = 16'h1ff;
			16'h854: y = 16'h1ff;
			16'h855: y = 16'h1ff;
			16'h856: y = 16'h1ff;
			16'h857: y = 16'h1ff;
			16'h858: y = 16'h1ff;
			16'h859: y = 16'h1ff;
			16'h85a: y = 16'h1ff;
			16'h85b: y = 16'h1ff;
			16'h85c: y = 16'h1ff;
			16'h85d: y = 16'h1ff;
			16'h85e: y = 16'h1ff;
			16'h85f: y = 16'h1ff;
			16'h860: y = 16'h1ff;
			16'h861: y = 16'h1ff;
			16'h862: y = 16'h1ff;
			16'h863: y = 16'h1ff;
			16'h864: y = 16'h1ff;
			16'h865: y = 16'h1ff;
			16'h866: y = 16'h1ff;
			16'h867: y = 16'h1ff;
			16'h868: y = 16'h1ff;
			16'h869: y = 16'h1ff;
			16'h86a: y = 16'h1ff;
			16'h86b: y = 16'h1ff;
			16'h86c: y = 16'h1ff;
			16'h86d: y = 16'h1ff;
			16'h86e: y = 16'h1ff;
			16'h86f: y = 16'h1ff;
			16'h870: y = 16'h1ff;
			16'h871: y = 16'h1ff;
			16'h872: y = 16'h1ff;
			16'h873: y = 16'h1ff;
			16'h874: y = 16'h1ff;
			16'h875: y = 16'h1ff;
			16'h876: y = 16'h1ff;
			16'h877: y = 16'h1ff;
			16'h878: y = 16'h1ff;
			16'h879: y = 16'h1ff;
			16'h87a: y = 16'h1ff;
			16'h87b: y = 16'h1ff;
			16'h87c: y = 16'h1ff;
			16'h87d: y = 16'h1ff;
			16'h87e: y = 16'h1ff;
			16'h87f: y = 16'h1ff;
			16'h880: y = 16'h1ff;
			16'h881: y = 16'h1ff;
			16'h882: y = 16'h1ff;
			16'h883: y = 16'h1ff;
			16'h884: y = 16'h1ff;
			16'h885: y = 16'h1ff;
			16'h886: y = 16'h1ff;
			16'h887: y = 16'h1ff;
			16'h888: y = 16'h1ff;
			16'h889: y = 16'h1ff;
			16'h88a: y = 16'h1ff;
			16'h88b: y = 16'h1ff;
			16'h88c: y = 16'h1ff;
			16'h88d: y = 16'h1ff;
			16'h88e: y = 16'h1ff;
			16'h88f: y = 16'h1ff;
			16'h890: y = 16'h1ff;
			16'h891: y = 16'h1ff;
			16'h892: y = 16'h1ff;
			16'h893: y = 16'h1ff;
			16'h894: y = 16'h1ff;
			16'h895: y = 16'h1ff;
			16'h896: y = 16'h1ff;
			16'h897: y = 16'h1ff;
			16'h898: y = 16'h1ff;
			16'h899: y = 16'h1ff;
			16'h89a: y = 16'h1ff;
			16'h89b: y = 16'h1ff;
			16'h89c: y = 16'h1ff;
			16'h89d: y = 16'h1ff;
			16'h89e: y = 16'h1ff;
			16'h89f: y = 16'h1ff;
			16'h8a0: y = 16'h1ff;
			16'h8a1: y = 16'h1ff;
			16'h8a2: y = 16'h1ff;
			16'h8a3: y = 16'h1ff;
			16'h8a4: y = 16'h1ff;
			16'h8a5: y = 16'h1ff;
			16'h8a6: y = 16'h1ff;
			16'h8a7: y = 16'h1ff;
			16'h8a8: y = 16'h1ff;
			16'h8a9: y = 16'h1ff;
			16'h8aa: y = 16'h1ff;
			16'h8ab: y = 16'h1ff;
			16'h8ac: y = 16'h1ff;
			16'h8ad: y = 16'h1ff;
			16'h8ae: y = 16'h1ff;
			16'h8af: y = 16'h1ff;
			16'h8b0: y = 16'h1ff;
			16'h8b1: y = 16'h1ff;
			16'h8b2: y = 16'h1ff;
			16'h8b3: y = 16'h1ff;
			16'h8b4: y = 16'h1ff;
			16'h8b5: y = 16'h1ff;
			16'h8b6: y = 16'h1ff;
			16'h8b7: y = 16'h1ff;
			16'h8b8: y = 16'h1ff;
			16'h8b9: y = 16'h1ff;
			16'h8ba: y = 16'h1ff;
			16'h8bb: y = 16'h1ff;
			16'h8bc: y = 16'h1ff;
			16'h8bd: y = 16'h1ff;
			16'h8be: y = 16'h1ff;
			16'h8bf: y = 16'h1ff;
			16'h8c0: y = 16'h1ff;
			16'h8c1: y = 16'h1ff;
			16'h8c2: y = 16'h1ff;
			16'h8c3: y = 16'h1ff;
			16'h8c4: y = 16'h1ff;
			16'h8c5: y = 16'h1ff;
			16'h8c6: y = 16'h1ff;
			16'h8c7: y = 16'h1ff;
			16'h8c8: y = 16'h1ff;
			16'h8c9: y = 16'h1ff;
			16'h8ca: y = 16'h1ff;
			16'h8cb: y = 16'h1ff;
			16'h8cc: y = 16'h1ff;
			16'h8cd: y = 16'h1ff;
			16'h8ce: y = 16'h1ff;
			16'h8cf: y = 16'h1ff;
			16'h8d0: y = 16'h1ff;
			16'h8d1: y = 16'h1ff;
			16'h8d2: y = 16'h1ff;
			16'h8d3: y = 16'h1ff;
			16'h8d4: y = 16'h1ff;
			16'h8d5: y = 16'h1ff;
			16'h8d6: y = 16'h1ff;
			16'h8d7: y = 16'h1ff;
			16'h8d8: y = 16'h1ff;
			16'h8d9: y = 16'h1ff;
			16'h8da: y = 16'h1ff;
			16'h8db: y = 16'h1ff;
			16'h8dc: y = 16'h1ff;
			16'h8dd: y = 16'h1ff;
			16'h8de: y = 16'h1ff;
			16'h8df: y = 16'h1ff;
			16'h8e0: y = 16'h1ff;
			16'h8e1: y = 16'h1ff;
			16'h8e2: y = 16'h1ff;
			16'h8e3: y = 16'h1ff;
			16'h8e4: y = 16'h1ff;
			16'h8e5: y = 16'h1ff;
			16'h8e6: y = 16'h1ff;
			16'h8e7: y = 16'h1ff;
			16'h8e8: y = 16'h1ff;
			16'h8e9: y = 16'h1ff;
			16'h8ea: y = 16'h1ff;
			16'h8eb: y = 16'h1ff;
			16'h8ec: y = 16'h1ff;
			16'h8ed: y = 16'h1ff;
			16'h8ee: y = 16'h1ff;
			16'h8ef: y = 16'h1ff;
			16'h8f0: y = 16'h1ff;
			16'h8f1: y = 16'h1ff;
			16'h8f2: y = 16'h1ff;
			16'h8f3: y = 16'h1ff;
			16'h8f4: y = 16'h1ff;
			16'h8f5: y = 16'h1ff;
			16'h8f6: y = 16'h1ff;
			16'h8f7: y = 16'h1ff;
			16'h8f8: y = 16'h1ff;
			16'h8f9: y = 16'h1ff;
			16'h8fa: y = 16'h1ff;
			16'h8fb: y = 16'h1ff;
			16'h8fc: y = 16'h1ff;
			16'h8fd: y = 16'h1ff;
			16'h8fe: y = 16'h1ff;
			16'h8ff: y = 16'h1ff;
			16'h900: y = 16'h1ff;
			16'h901: y = 16'h1ff;
			16'h902: y = 16'h1ff;
			16'h903: y = 16'h1ff;
			16'h904: y = 16'h1ff;
			16'h905: y = 16'h1ff;
			16'h906: y = 16'h1ff;
			16'h907: y = 16'h1ff;
			16'h908: y = 16'h1ff;
			16'h909: y = 16'h1ff;
			16'h90a: y = 16'h1ff;
			16'h90b: y = 16'h1ff;
			16'h90c: y = 16'h1ff;
			16'h90d: y = 16'h1ff;
			16'h90e: y = 16'h1ff;
			16'h90f: y = 16'h1ff;
			16'h910: y = 16'h1ff;
			16'h911: y = 16'h1ff;
			16'h912: y = 16'h1ff;
			16'h913: y = 16'h1ff;
			16'h914: y = 16'h1ff;
			16'h915: y = 16'h1ff;
			16'h916: y = 16'h1ff;
			16'h917: y = 16'h1ff;
			16'h918: y = 16'h1ff;
			16'h919: y = 16'h1ff;
			16'h91a: y = 16'h1ff;
			16'h91b: y = 16'h1ff;
			16'h91c: y = 16'h1ff;
			16'h91d: y = 16'h1ff;
			16'h91e: y = 16'h1ff;
			16'h91f: y = 16'h1ff;
			16'h920: y = 16'h1ff;
			16'h921: y = 16'h1ff;
			16'h922: y = 16'h1ff;
			16'h923: y = 16'h1ff;
			16'h924: y = 16'h1ff;
			16'h925: y = 16'h1ff;
			16'h926: y = 16'h1ff;
			16'h927: y = 16'h1ff;
			16'h928: y = 16'h1ff;
			16'h929: y = 16'h1ff;
			16'h92a: y = 16'h1ff;
			16'h92b: y = 16'h1ff;
			16'h92c: y = 16'h1ff;
			16'h92d: y = 16'h1ff;
			16'h92e: y = 16'h1ff;
			16'h92f: y = 16'h1ff;
			16'h930: y = 16'h1ff;
			16'h931: y = 16'h1ff;
			16'h932: y = 16'h1ff;
			16'h933: y = 16'h1ff;
			16'h934: y = 16'h1ff;
			16'h935: y = 16'h1ff;
			16'h936: y = 16'h1ff;
			16'h937: y = 16'h1ff;
			16'h938: y = 16'h1ff;
			16'h939: y = 16'h1ff;
			16'h93a: y = 16'h1ff;
			16'h93b: y = 16'h1ff;
			16'h93c: y = 16'h1ff;
			16'h93d: y = 16'h1ff;
			16'h93e: y = 16'h1ff;
			16'h93f: y = 16'h1ff;
			16'h940: y = 16'h1ff;
			16'h941: y = 16'h1ff;
			16'h942: y = 16'h1ff;
			16'h943: y = 16'h1ff;
			16'h944: y = 16'h1ff;
			16'h945: y = 16'h1ff;
			16'h946: y = 16'h1ff;
			16'h947: y = 16'h1ff;
			16'h948: y = 16'h1ff;
			16'h949: y = 16'h1ff;
			16'h94a: y = 16'h1ff;
			16'h94b: y = 16'h1ff;
			16'h94c: y = 16'h1ff;
			16'h94d: y = 16'h1ff;
			16'h94e: y = 16'h1ff;
			16'h94f: y = 16'h1ff;
			16'h950: y = 16'h1ff;
			16'h951: y = 16'h1ff;
			16'h952: y = 16'h1ff;
			16'h953: y = 16'h1ff;
			16'h954: y = 16'h1ff;
			16'h955: y = 16'h1ff;
			16'h956: y = 16'h1ff;
			16'h957: y = 16'h1ff;
			16'h958: y = 16'h1ff;
			16'h959: y = 16'h1ff;
			16'h95a: y = 16'h1ff;
			16'h95b: y = 16'h1ff;
			16'h95c: y = 16'h1ff;
			16'h95d: y = 16'h1ff;
			16'h95e: y = 16'h1ff;
			16'h95f: y = 16'h1ff;
			16'h960: y = 16'h1ff;
			16'h961: y = 16'h1ff;
			16'h962: y = 16'h1ff;
			16'h963: y = 16'h1ff;
			16'h964: y = 16'h1ff;
			16'h965: y = 16'h1ff;
			16'h966: y = 16'h1ff;
			16'h967: y = 16'h1ff;
			16'h968: y = 16'h1ff;
			16'h969: y = 16'h1ff;
			16'h96a: y = 16'h1ff;
			16'h96b: y = 16'h1ff;
			16'h96c: y = 16'h1ff;
			16'h96d: y = 16'h1ff;
			16'h96e: y = 16'h1ff;
			16'h96f: y = 16'h1ff;
			16'h970: y = 16'h1ff;
			16'h971: y = 16'h1ff;
			16'h972: y = 16'h1ff;
			16'h973: y = 16'h1ff;
			16'h974: y = 16'h1ff;
			16'h975: y = 16'h1ff;
			16'h976: y = 16'h1ff;
			16'h977: y = 16'h1ff;
			16'h978: y = 16'h1ff;
			16'h979: y = 16'h1ff;
			16'h97a: y = 16'h1ff;
			16'h97b: y = 16'h1ff;
			16'h97c: y = 16'h1ff;
			16'h97d: y = 16'h1ff;
			16'h97e: y = 16'h1ff;
			16'h97f: y = 16'h1ff;
			16'h980: y = 16'h1ff;
			16'h981: y = 16'h1ff;
			16'h982: y = 16'h1ff;
			16'h983: y = 16'h1ff;
			16'h984: y = 16'h1ff;
			16'h985: y = 16'h1ff;
			16'h986: y = 16'h1ff;
			16'h987: y = 16'h1ff;
			16'h988: y = 16'h1ff;
			16'h989: y = 16'h1ff;
			16'h98a: y = 16'h1ff;
			16'h98b: y = 16'h1ff;
			16'h98c: y = 16'h1ff;
			16'h98d: y = 16'h1ff;
			16'h98e: y = 16'h1ff;
			16'h98f: y = 16'h1ff;
			16'h990: y = 16'h1ff;
			16'h991: y = 16'h1ff;
			16'h992: y = 16'h1ff;
			16'h993: y = 16'h1ff;
			16'h994: y = 16'h1ff;
			16'h995: y = 16'h1ff;
			16'h996: y = 16'h1ff;
			16'h997: y = 16'h1ff;
			16'h998: y = 16'h1ff;
			16'h999: y = 16'h1ff;
			16'h99a: y = 16'h1ff;
			16'h99b: y = 16'h1ff;
			16'h99c: y = 16'h1ff;
			16'h99d: y = 16'h1ff;
			16'h99e: y = 16'h1ff;
			16'h99f: y = 16'h1ff;
			16'h9a0: y = 16'h1ff;
			16'h9a1: y = 16'h1ff;
			16'h9a2: y = 16'h1ff;
			16'h9a3: y = 16'h1ff;
			16'h9a4: y = 16'h1ff;
			16'h9a5: y = 16'h1ff;
			16'h9a6: y = 16'h1ff;
			16'h9a7: y = 16'h1ff;
			16'h9a8: y = 16'h1ff;
			16'h9a9: y = 16'h1ff;
			16'h9aa: y = 16'h1ff;
			16'h9ab: y = 16'h1ff;
			16'h9ac: y = 16'h1ff;
			16'h9ad: y = 16'h1ff;
			16'h9ae: y = 16'h1ff;
			16'h9af: y = 16'h1ff;
			16'h9b0: y = 16'h1ff;
			16'h9b1: y = 16'h1ff;
			16'h9b2: y = 16'h1ff;
			16'h9b3: y = 16'h1ff;
			16'h9b4: y = 16'h1ff;
			16'h9b5: y = 16'h1ff;
			16'h9b6: y = 16'h1ff;
			16'h9b7: y = 16'h1ff;
			16'h9b8: y = 16'h1ff;
			16'h9b9: y = 16'h1ff;
			16'h9ba: y = 16'h1ff;
			16'h9bb: y = 16'h1ff;
			16'h9bc: y = 16'h1ff;
			16'h9bd: y = 16'h1ff;
			16'h9be: y = 16'h1ff;
			16'h9bf: y = 16'h1ff;
			16'h9c0: y = 16'h1ff;
			16'h9c1: y = 16'h1ff;
			16'h9c2: y = 16'h1ff;
			16'h9c3: y = 16'h1ff;
			16'h9c4: y = 16'h1ff;
			16'h9c5: y = 16'h1ff;
			16'h9c6: y = 16'h1ff;
			16'h9c7: y = 16'h1ff;
			16'h9c8: y = 16'h1ff;
			16'h9c9: y = 16'h1ff;
			16'h9ca: y = 16'h1ff;
			16'h9cb: y = 16'h1ff;
			16'h9cc: y = 16'h1ff;
			16'h9cd: y = 16'h1ff;
			16'h9ce: y = 16'h1ff;
			16'h9cf: y = 16'h1ff;
			16'h9d0: y = 16'h1ff;
			16'h9d1: y = 16'h1ff;
			16'h9d2: y = 16'h1ff;
			16'h9d3: y = 16'h1ff;
			16'h9d4: y = 16'h1ff;
			16'h9d5: y = 16'h1ff;
			16'h9d6: y = 16'h1ff;
			16'h9d7: y = 16'h1ff;
			16'h9d8: y = 16'h1ff;
			16'h9d9: y = 16'h1ff;
			16'h9da: y = 16'h1ff;
			16'h9db: y = 16'h1ff;
			16'h9dc: y = 16'h1ff;
			16'h9dd: y = 16'h1ff;
			16'h9de: y = 16'h1ff;
			16'h9df: y = 16'h1ff;
			16'h9e0: y = 16'h1ff;
			16'h9e1: y = 16'h1ff;
			16'h9e2: y = 16'h1ff;
			16'h9e3: y = 16'h1ff;
			16'h9e4: y = 16'h1ff;
			16'h9e5: y = 16'h1ff;
			16'h9e6: y = 16'h1ff;
			16'h9e7: y = 16'h1ff;
			16'h9e8: y = 16'h1ff;
			16'h9e9: y = 16'h1ff;
			16'h9ea: y = 16'h1ff;
			16'h9eb: y = 16'h1ff;
			16'h9ec: y = 16'h1ff;
			16'h9ed: y = 16'h1ff;
			16'h9ee: y = 16'h1ff;
			16'h9ef: y = 16'h1ff;
			16'h9f0: y = 16'h1ff;
			16'h9f1: y = 16'h1ff;
			16'h9f2: y = 16'h1ff;
			16'h9f3: y = 16'h1ff;
			16'h9f4: y = 16'h1ff;
			16'h9f5: y = 16'h1ff;
			16'h9f6: y = 16'h1ff;
			16'h9f7: y = 16'h1ff;
			16'h9f8: y = 16'h1ff;
			16'h9f9: y = 16'h1ff;
			16'h9fa: y = 16'h1ff;
			16'h9fb: y = 16'h1ff;
			16'h9fc: y = 16'h1ff;
			16'h9fd: y = 16'h1ff;
			16'h9fe: y = 16'h1ff;
			16'h9ff: y = 16'h1ff;
			16'ha00: y = 16'h1ff;
			16'ha01: y = 16'h1ff;
			16'ha02: y = 16'h1ff;
			16'ha03: y = 16'h1ff;
			16'ha04: y = 16'h1ff;
			16'ha05: y = 16'h1ff;
			16'ha06: y = 16'h1ff;
			16'ha07: y = 16'h1ff;
			16'ha08: y = 16'h1ff;
			16'ha09: y = 16'h1ff;
			16'ha0a: y = 16'h1ff;
			16'ha0b: y = 16'h1ff;
			16'ha0c: y = 16'h1ff;
			16'ha0d: y = 16'h1ff;
			16'ha0e: y = 16'h1ff;
			16'ha0f: y = 16'h1ff;
			16'ha10: y = 16'h1ff;
			16'ha11: y = 16'h1ff;
			16'ha12: y = 16'h1ff;
			16'ha13: y = 16'h1ff;
			16'ha14: y = 16'h1ff;
			16'ha15: y = 16'h1ff;
			16'ha16: y = 16'h1ff;
			16'ha17: y = 16'h1ff;
			16'ha18: y = 16'h1ff;
			16'ha19: y = 16'h1ff;
			16'ha1a: y = 16'h1ff;
			16'ha1b: y = 16'h1ff;
			16'ha1c: y = 16'h1ff;
			16'ha1d: y = 16'h1ff;
			16'ha1e: y = 16'h1ff;
			16'ha1f: y = 16'h1ff;
			16'ha20: y = 16'h1ff;
			16'ha21: y = 16'h1ff;
			16'ha22: y = 16'h1ff;
			16'ha23: y = 16'h1ff;
			16'ha24: y = 16'h1ff;
			16'ha25: y = 16'h1ff;
			16'ha26: y = 16'h1ff;
			16'ha27: y = 16'h1ff;
			16'ha28: y = 16'h1ff;
			16'ha29: y = 16'h1ff;
			16'ha2a: y = 16'h1ff;
			16'ha2b: y = 16'h1ff;
			16'ha2c: y = 16'h1ff;
			16'ha2d: y = 16'h1ff;
			16'ha2e: y = 16'h1ff;
			16'ha2f: y = 16'h1ff;
			16'ha30: y = 16'h1ff;
			16'ha31: y = 16'h1ff;
			16'ha32: y = 16'h1ff;
			16'ha33: y = 16'h1ff;
			16'ha34: y = 16'h1ff;
			16'ha35: y = 16'h1ff;
			16'ha36: y = 16'h1ff;
			16'ha37: y = 16'h1ff;
			16'ha38: y = 16'h1ff;
			16'ha39: y = 16'h1ff;
			16'ha3a: y = 16'h1ff;
			16'ha3b: y = 16'h1ff;
			16'ha3c: y = 16'h1ff;
			16'ha3d: y = 16'h1ff;
			16'ha3e: y = 16'h1ff;
			16'ha3f: y = 16'h1ff;
			16'ha40: y = 16'h1ff;
			16'ha41: y = 16'h1ff;
			16'ha42: y = 16'h1ff;
			16'ha43: y = 16'h1ff;
			16'ha44: y = 16'h1ff;
			16'ha45: y = 16'h1ff;
			16'ha46: y = 16'h1ff;
			16'ha47: y = 16'h1ff;
			16'ha48: y = 16'h1ff;
			16'ha49: y = 16'h1ff;
			16'ha4a: y = 16'h1ff;
			16'ha4b: y = 16'h1ff;
			16'ha4c: y = 16'h1ff;
			16'ha4d: y = 16'h1ff;
			16'ha4e: y = 16'h1ff;
			16'ha4f: y = 16'h1ff;
			16'ha50: y = 16'h1ff;
			16'ha51: y = 16'h1ff;
			16'ha52: y = 16'h1ff;
			16'ha53: y = 16'h1ff;
			16'ha54: y = 16'h1ff;
			16'ha55: y = 16'h1ff;
			16'ha56: y = 16'h1ff;
			16'ha57: y = 16'h1ff;
			16'ha58: y = 16'h1ff;
			16'ha59: y = 16'h1ff;
			16'ha5a: y = 16'h1ff;
			16'ha5b: y = 16'h1ff;
			16'ha5c: y = 16'h1ff;
			16'ha5d: y = 16'h1ff;
			16'ha5e: y = 16'h1ff;
			16'ha5f: y = 16'h1ff;
			16'ha60: y = 16'h1ff;
			16'ha61: y = 16'h1ff;
			16'ha62: y = 16'h1ff;
			16'ha63: y = 16'h1ff;
			16'ha64: y = 16'h1ff;
			16'ha65: y = 16'h1ff;
			16'ha66: y = 16'h1ff;
			16'ha67: y = 16'h1ff;
			16'ha68: y = 16'h1ff;
			16'ha69: y = 16'h1ff;
			16'ha6a: y = 16'h1ff;
			16'ha6b: y = 16'h1ff;
			16'ha6c: y = 16'h1ff;
			16'ha6d: y = 16'h1ff;
			16'ha6e: y = 16'h1ff;
			16'ha6f: y = 16'h1ff;
			16'ha70: y = 16'h1ff;
			16'ha71: y = 16'h1ff;
			16'ha72: y = 16'h1ff;
			16'ha73: y = 16'h1ff;
			16'ha74: y = 16'h1ff;
			16'ha75: y = 16'h1ff;
			16'ha76: y = 16'h1ff;
			16'ha77: y = 16'h1ff;
			16'ha78: y = 16'h1ff;
			16'ha79: y = 16'h1ff;
			16'ha7a: y = 16'h1ff;
			16'ha7b: y = 16'h1ff;
			16'ha7c: y = 16'h1ff;
			16'ha7d: y = 16'h1ff;
			16'ha7e: y = 16'h1ff;
			16'ha7f: y = 16'h1ff;
			16'ha80: y = 16'h1ff;
			16'ha81: y = 16'h1ff;
			16'ha82: y = 16'h1ff;
			16'ha83: y = 16'h1ff;
			16'ha84: y = 16'h1ff;
			16'ha85: y = 16'h1ff;
			16'ha86: y = 16'h1ff;
			16'ha87: y = 16'h1ff;
			16'ha88: y = 16'h1ff;
			16'ha89: y = 16'h1ff;
			16'ha8a: y = 16'h1ff;
			16'ha8b: y = 16'h1ff;
			16'ha8c: y = 16'h1ff;
			16'ha8d: y = 16'h1ff;
			16'ha8e: y = 16'h1ff;
			16'ha8f: y = 16'h1ff;
			16'ha90: y = 16'h1ff;
			16'ha91: y = 16'h1ff;
			16'ha92: y = 16'h1ff;
			16'ha93: y = 16'h1ff;
			16'ha94: y = 16'h1ff;
			16'ha95: y = 16'h1ff;
			16'ha96: y = 16'h1ff;
			16'ha97: y = 16'h1ff;
			16'ha98: y = 16'h1ff;
			16'ha99: y = 16'h1ff;
			16'ha9a: y = 16'h1ff;
			16'ha9b: y = 16'h1ff;
			16'ha9c: y = 16'h1ff;
			16'ha9d: y = 16'h1ff;
			16'ha9e: y = 16'h1ff;
			16'ha9f: y = 16'h1ff;
			16'haa0: y = 16'h1ff;
			16'haa1: y = 16'h1ff;
			16'haa2: y = 16'h1ff;
			16'haa3: y = 16'h1ff;
			16'haa4: y = 16'h1ff;
			16'haa5: y = 16'h1ff;
			16'haa6: y = 16'h1ff;
			16'haa7: y = 16'h1ff;
			16'haa8: y = 16'h1ff;
			16'haa9: y = 16'h1ff;
			16'haaa: y = 16'h1ff;
			16'haab: y = 16'h1ff;
			16'haac: y = 16'h1ff;
			16'haad: y = 16'h1ff;
			16'haae: y = 16'h1ff;
			16'haaf: y = 16'h1ff;
			16'hab0: y = 16'h1ff;
			16'hab1: y = 16'h1ff;
			16'hab2: y = 16'h1ff;
			16'hab3: y = 16'h1ff;
			16'hab4: y = 16'h1ff;
			16'hab5: y = 16'h1ff;
			16'hab6: y = 16'h1ff;
			16'hab7: y = 16'h1ff;
			16'hab8: y = 16'h1ff;
			16'hab9: y = 16'h1ff;
			16'haba: y = 16'h1ff;
			16'habb: y = 16'h1ff;
			16'habc: y = 16'h1ff;
			16'habd: y = 16'h1ff;
			16'habe: y = 16'h1ff;
			16'habf: y = 16'h1ff;
			16'hac0: y = 16'h1ff;
			16'hac1: y = 16'h1ff;
			16'hac2: y = 16'h1ff;
			16'hac3: y = 16'h1ff;
			16'hac4: y = 16'h1ff;
			16'hac5: y = 16'h1ff;
			16'hac6: y = 16'h1ff;
			16'hac7: y = 16'h1ff;
			16'hac8: y = 16'h1ff;
			16'hac9: y = 16'h1ff;
			16'haca: y = 16'h1ff;
			16'hacb: y = 16'h1ff;
			16'hacc: y = 16'h1ff;
			16'hacd: y = 16'h1ff;
			16'hace: y = 16'h1ff;
			16'hacf: y = 16'h1ff;
			16'had0: y = 16'h1ff;
			16'had1: y = 16'h1ff;
			16'had2: y = 16'h1ff;
			16'had3: y = 16'h1ff;
			16'had4: y = 16'h1ff;
			16'had5: y = 16'h1ff;
			16'had6: y = 16'h1ff;
			16'had7: y = 16'h1ff;
			16'had8: y = 16'h1ff;
			16'had9: y = 16'h1ff;
			16'hada: y = 16'h1ff;
			16'hadb: y = 16'h1ff;
			16'hadc: y = 16'h1ff;
			16'hadd: y = 16'h1ff;
			16'hade: y = 16'h1ff;
			16'hadf: y = 16'h1ff;
			16'hae0: y = 16'h1ff;
			16'hae1: y = 16'h1ff;
			16'hae2: y = 16'h1ff;
			16'hae3: y = 16'h1ff;
			16'hae4: y = 16'h1ff;
			16'hae5: y = 16'h1ff;
			16'hae6: y = 16'h1ff;
			16'hae7: y = 16'h1ff;
			16'hae8: y = 16'h1ff;
			16'hae9: y = 16'h1ff;
			16'haea: y = 16'h1ff;
			16'haeb: y = 16'h1ff;
			16'haec: y = 16'h1ff;
			16'haed: y = 16'h1ff;
			16'haee: y = 16'h1ff;
			16'haef: y = 16'h1ff;
			16'haf0: y = 16'h1ff;
			16'haf1: y = 16'h1ff;
			16'haf2: y = 16'h1ff;
			16'haf3: y = 16'h1ff;
			16'haf4: y = 16'h1ff;
			16'haf5: y = 16'h1ff;
			16'haf6: y = 16'h1ff;
			16'haf7: y = 16'h1ff;
			16'haf8: y = 16'h1ff;
			16'haf9: y = 16'h1ff;
			16'hafa: y = 16'h1ff;
			16'hafb: y = 16'h1ff;
			16'hafc: y = 16'h1ff;
			16'hafd: y = 16'h1ff;
			16'hafe: y = 16'h1ff;
			16'haff: y = 16'h1ff;
			16'hb00: y = 16'h1ff;
			16'hb01: y = 16'h1ff;
			16'hb02: y = 16'h1ff;
			16'hb03: y = 16'h1ff;
			16'hb04: y = 16'h1ff;
			16'hb05: y = 16'h1ff;
			16'hb06: y = 16'h1ff;
			16'hb07: y = 16'h1ff;
			16'hb08: y = 16'h1ff;
			16'hb09: y = 16'h1ff;
			16'hb0a: y = 16'h1ff;
			16'hb0b: y = 16'h1ff;
			16'hb0c: y = 16'h1ff;
			16'hb0d: y = 16'h1ff;
			16'hb0e: y = 16'h1ff;
			16'hb0f: y = 16'h1ff;
			16'hb10: y = 16'h1ff;
			16'hb11: y = 16'h1ff;
			16'hb12: y = 16'h1ff;
			16'hb13: y = 16'h1ff;
			16'hb14: y = 16'h1ff;
			16'hb15: y = 16'h1ff;
			16'hb16: y = 16'h1ff;
			16'hb17: y = 16'h1ff;
			16'hb18: y = 16'h1ff;
			16'hb19: y = 16'h1ff;
			16'hb1a: y = 16'h1ff;
			16'hb1b: y = 16'h1ff;
			16'hb1c: y = 16'h1ff;
			16'hb1d: y = 16'h1ff;
			16'hb1e: y = 16'h1ff;
			16'hb1f: y = 16'h1ff;
			16'hb20: y = 16'h1ff;
			16'hb21: y = 16'h1ff;
			16'hb22: y = 16'h1ff;
			16'hb23: y = 16'h1ff;
			16'hb24: y = 16'h1ff;
			16'hb25: y = 16'h1ff;
			16'hb26: y = 16'h1ff;
			16'hb27: y = 16'h1ff;
			16'hb28: y = 16'h1ff;
			16'hb29: y = 16'h1ff;
			16'hb2a: y = 16'h1ff;
			16'hb2b: y = 16'h1ff;
			16'hb2c: y = 16'h1ff;
			16'hb2d: y = 16'h1ff;
			16'hb2e: y = 16'h1ff;
			16'hb2f: y = 16'h1ff;
			16'hb30: y = 16'h1ff;
			16'hb31: y = 16'h1ff;
			16'hb32: y = 16'h1ff;
			16'hb33: y = 16'h1ff;
			16'hb34: y = 16'h1ff;
			16'hb35: y = 16'h1ff;
			16'hb36: y = 16'h1ff;
			16'hb37: y = 16'h1ff;
			16'hb38: y = 16'h1ff;
			16'hb39: y = 16'h1ff;
			16'hb3a: y = 16'h1ff;
			16'hb3b: y = 16'h1ff;
			16'hb3c: y = 16'h1ff;
			16'hb3d: y = 16'h1ff;
			16'hb3e: y = 16'h1ff;
			16'hb3f: y = 16'h1ff;
			16'hb40: y = 16'h1ff;
			16'hb41: y = 16'h1ff;
			16'hb42: y = 16'h1ff;
			16'hb43: y = 16'h1ff;
			16'hb44: y = 16'h1ff;
			16'hb45: y = 16'h1ff;
			16'hb46: y = 16'h1ff;
			16'hb47: y = 16'h1ff;
			16'hb48: y = 16'h1ff;
			16'hb49: y = 16'h1ff;
			16'hb4a: y = 16'h1ff;
			16'hb4b: y = 16'h1ff;
			16'hb4c: y = 16'h1ff;
			16'hb4d: y = 16'h1ff;
			16'hb4e: y = 16'h1ff;
			16'hb4f: y = 16'h1ff;
			16'hb50: y = 16'h1ff;
			16'hb51: y = 16'h1ff;
			16'hb52: y = 16'h1ff;
			16'hb53: y = 16'h1ff;
			16'hb54: y = 16'h1ff;
			16'hb55: y = 16'h1ff;
			16'hb56: y = 16'h1ff;
			16'hb57: y = 16'h1ff;
			16'hb58: y = 16'h1ff;
			16'hb59: y = 16'h1ff;
			16'hb5a: y = 16'h1ff;
			16'hb5b: y = 16'h1ff;
			16'hb5c: y = 16'h1ff;
			16'hb5d: y = 16'h1ff;
			16'hb5e: y = 16'h1ff;
			16'hb5f: y = 16'h1ff;
			16'hb60: y = 16'h1ff;
			16'hb61: y = 16'h1ff;
			16'hb62: y = 16'h1ff;
			16'hb63: y = 16'h1ff;
			16'hb64: y = 16'h1ff;
			16'hb65: y = 16'h1ff;
			16'hb66: y = 16'h1ff;
			16'hb67: y = 16'h1ff;
			16'hb68: y = 16'h1ff;
			16'hb69: y = 16'h1ff;
			16'hb6a: y = 16'h1ff;
			16'hb6b: y = 16'h1ff;
			16'hb6c: y = 16'h1ff;
			16'hb6d: y = 16'h1ff;
			16'hb6e: y = 16'h1ff;
			16'hb6f: y = 16'h1ff;
			16'hb70: y = 16'h1ff;
			16'hb71: y = 16'h1ff;
			16'hb72: y = 16'h1ff;
			16'hb73: y = 16'h1ff;
			16'hb74: y = 16'h1ff;
			16'hb75: y = 16'h1ff;
			16'hb76: y = 16'h1ff;
			16'hb77: y = 16'h1ff;
			16'hb78: y = 16'h1ff;
			16'hb79: y = 16'h1ff;
			16'hb7a: y = 16'h1ff;
			16'hb7b: y = 16'h1ff;
			16'hb7c: y = 16'h1ff;
			16'hb7d: y = 16'h1ff;
			16'hb7e: y = 16'h1ff;
			16'hb7f: y = 16'h1ff;
			16'hb80: y = 16'h1ff;
			16'hb81: y = 16'h1ff;
			16'hb82: y = 16'h1ff;
			16'hb83: y = 16'h1ff;
			16'hb84: y = 16'h1ff;
			16'hb85: y = 16'h1ff;
			16'hb86: y = 16'h1ff;
			16'hb87: y = 16'h1ff;
			16'hb88: y = 16'h1ff;
			16'hb89: y = 16'h1ff;
			16'hb8a: y = 16'h1ff;
			16'hb8b: y = 16'h1ff;
			16'hb8c: y = 16'h1ff;
			16'hb8d: y = 16'h1ff;
			16'hb8e: y = 16'h1ff;
			16'hb8f: y = 16'h1ff;
			16'hb90: y = 16'h1ff;
			16'hb91: y = 16'h1ff;
			16'hb92: y = 16'h1ff;
			16'hb93: y = 16'h1ff;
			16'hb94: y = 16'h1ff;
			16'hb95: y = 16'h1ff;
			16'hb96: y = 16'h1ff;
			16'hb97: y = 16'h1ff;
			16'hb98: y = 16'h1ff;
			16'hb99: y = 16'h1ff;
			16'hb9a: y = 16'h1ff;
			16'hb9b: y = 16'h1ff;
			16'hb9c: y = 16'h1ff;
			16'hb9d: y = 16'h1ff;
			16'hb9e: y = 16'h1ff;
			16'hb9f: y = 16'h1ff;
			16'hba0: y = 16'h1ff;
			16'hba1: y = 16'h1ff;
			16'hba2: y = 16'h1ff;
			16'hba3: y = 16'h1ff;
			16'hba4: y = 16'h1ff;
			16'hba5: y = 16'h1ff;
			16'hba6: y = 16'h1ff;
			16'hba7: y = 16'h1ff;
			16'hba8: y = 16'h1ff;
			16'hba9: y = 16'h1ff;
			16'hbaa: y = 16'h1ff;
			16'hbab: y = 16'h1ff;
			16'hbac: y = 16'h1ff;
			16'hbad: y = 16'h1ff;
			16'hbae: y = 16'h1ff;
			16'hbaf: y = 16'h1ff;
			16'hbb0: y = 16'h1ff;
			16'hbb1: y = 16'h1ff;
			16'hbb2: y = 16'h1ff;
			16'hbb3: y = 16'h1ff;
			16'hbb4: y = 16'h1ff;
			16'hbb5: y = 16'h1ff;
			16'hbb6: y = 16'h1ff;
			16'hbb7: y = 16'h1ff;
			16'hbb8: y = 16'h1ff;
			16'hbb9: y = 16'h1ff;
			16'hbba: y = 16'h1ff;
			16'hbbb: y = 16'h1ff;
			16'hbbc: y = 16'h1ff;
			16'hbbd: y = 16'h1ff;
			16'hbbe: y = 16'h1ff;
			16'hbbf: y = 16'h1ff;
			16'hbc0: y = 16'h1ff;
			16'hbc1: y = 16'h1ff;
			16'hbc2: y = 16'h1ff;
			16'hbc3: y = 16'h1ff;
			16'hbc4: y = 16'h1ff;
			16'hbc5: y = 16'h1ff;
			16'hbc6: y = 16'h1ff;
			16'hbc7: y = 16'h1ff;
			16'hbc8: y = 16'h1ff;
			16'hbc9: y = 16'h1ff;
			16'hbca: y = 16'h1ff;
			16'hbcb: y = 16'h1ff;
			16'hbcc: y = 16'h1ff;
			16'hbcd: y = 16'h1ff;
			16'hbce: y = 16'h1ff;
			16'hbcf: y = 16'h1ff;
			16'hbd0: y = 16'h1ff;
			16'hbd1: y = 16'h1ff;
			16'hbd2: y = 16'h1ff;
			16'hbd3: y = 16'h1ff;
			16'hbd4: y = 16'h1ff;
			16'hbd5: y = 16'h1ff;
			16'hbd6: y = 16'h1ff;
			16'hbd7: y = 16'h1ff;
			16'hbd8: y = 16'h1ff;
			16'hbd9: y = 16'h1ff;
			16'hbda: y = 16'h1ff;
			16'hbdb: y = 16'h1ff;
			16'hbdc: y = 16'h1ff;
			16'hbdd: y = 16'h1ff;
			16'hbde: y = 16'h1ff;
			16'hbdf: y = 16'h1ff;
			16'hbe0: y = 16'h1ff;
			16'hbe1: y = 16'h1ff;
			16'hbe2: y = 16'h1ff;
			16'hbe3: y = 16'h1ff;
			16'hbe4: y = 16'h1ff;
			16'hbe5: y = 16'h1ff;
			16'hbe6: y = 16'h1ff;
			16'hbe7: y = 16'h1ff;
			16'hbe8: y = 16'h1ff;
			16'hbe9: y = 16'h1ff;
			16'hbea: y = 16'h1ff;
			16'hbeb: y = 16'h1ff;
			16'hbec: y = 16'h1ff;
			16'hbed: y = 16'h1ff;
			16'hbee: y = 16'h1ff;
			16'hbef: y = 16'h1ff;
			16'hbf0: y = 16'h1ff;
			16'hbf1: y = 16'h1ff;
			16'hbf2: y = 16'h1ff;
			16'hbf3: y = 16'h1ff;
			16'hbf4: y = 16'h1ff;
			16'hbf5: y = 16'h1ff;
			16'hbf6: y = 16'h1ff;
			16'hbf7: y = 16'h1ff;
			16'hbf8: y = 16'h1ff;
			16'hbf9: y = 16'h1ff;
			16'hbfa: y = 16'h1ff;
			16'hbfb: y = 16'h1ff;
			16'hbfc: y = 16'h1ff;
			16'hbfd: y = 16'h1ff;
			16'hbfe: y = 16'h1ff;
			16'hbff: y = 16'h1ff;
			16'hc00: y = 16'h1ff;
			16'hc01: y = 16'h1ff;
			16'hc02: y = 16'h1ff;
			16'hc03: y = 16'h1ff;
			16'hc04: y = 16'h1ff;
			16'hc05: y = 16'h1ff;
			16'hc06: y = 16'h1ff;
			16'hc07: y = 16'h1ff;
			16'hc08: y = 16'h1ff;
			16'hc09: y = 16'h1ff;
			16'hc0a: y = 16'h1ff;
			16'hc0b: y = 16'h1ff;
			16'hc0c: y = 16'h1ff;
			16'hc0d: y = 16'h1ff;
			16'hc0e: y = 16'h1ff;
			16'hc0f: y = 16'h1ff;
			16'hc10: y = 16'h1ff;
			16'hc11: y = 16'h1ff;
			16'hc12: y = 16'h1ff;
			16'hc13: y = 16'h1ff;
			16'hc14: y = 16'h1ff;
			16'hc15: y = 16'h1ff;
			16'hc16: y = 16'h1ff;
			16'hc17: y = 16'h1ff;
			16'hc18: y = 16'h1ff;
			16'hc19: y = 16'h1ff;
			16'hc1a: y = 16'h1ff;
			16'hc1b: y = 16'h1ff;
			16'hc1c: y = 16'h1ff;
			16'hc1d: y = 16'h1ff;
			16'hc1e: y = 16'h1ff;
			16'hc1f: y = 16'h1ff;
			16'hc20: y = 16'h1ff;
			16'hc21: y = 16'h1ff;
			16'hc22: y = 16'h1ff;
			16'hc23: y = 16'h1ff;
			16'hc24: y = 16'h1ff;
			16'hc25: y = 16'h1ff;
			16'hc26: y = 16'h1ff;
			16'hc27: y = 16'h1ff;
			16'hc28: y = 16'h1ff;
			16'hc29: y = 16'h1ff;
			16'hc2a: y = 16'h1ff;
			16'hc2b: y = 16'h1ff;
			16'hc2c: y = 16'h1ff;
			16'hc2d: y = 16'h1ff;
			16'hc2e: y = 16'h1ff;
			16'hc2f: y = 16'h1ff;
			16'hc30: y = 16'h1ff;
			16'hc31: y = 16'h1ff;
			16'hc32: y = 16'h1ff;
			16'hc33: y = 16'h1ff;
			16'hc34: y = 16'h1ff;
			16'hc35: y = 16'h1ff;
			16'hc36: y = 16'h1ff;
			16'hc37: y = 16'h1ff;
			16'hc38: y = 16'h1ff;
			16'hc39: y = 16'h1ff;
			16'hc3a: y = 16'h1ff;
			16'hc3b: y = 16'h1ff;
			16'hc3c: y = 16'h1ff;
			16'hc3d: y = 16'h1ff;
			16'hc3e: y = 16'h1ff;
			16'hc3f: y = 16'h1ff;
			16'hc40: y = 16'h1ff;
			16'hc41: y = 16'h1ff;
			16'hc42: y = 16'h1ff;
			16'hc43: y = 16'h1ff;
			16'hc44: y = 16'h1ff;
			16'hc45: y = 16'h1ff;
			16'hc46: y = 16'h1ff;
			16'hc47: y = 16'h1ff;
			16'hc48: y = 16'h1ff;
			16'hc49: y = 16'h1ff;
			16'hc4a: y = 16'h1ff;
			16'hc4b: y = 16'h1ff;
			16'hc4c: y = 16'h1ff;
			16'hc4d: y = 16'h1ff;
			16'hc4e: y = 16'h1ff;
			16'hc4f: y = 16'h1ff;
			16'hc50: y = 16'h1ff;
			16'hc51: y = 16'h1ff;
			16'hc52: y = 16'h1ff;
			16'hc53: y = 16'h1ff;
			16'hc54: y = 16'h1ff;
			16'hc55: y = 16'h1ff;
			16'hc56: y = 16'h1ff;
			16'hc57: y = 16'h1ff;
			16'hc58: y = 16'h1ff;
			16'hc59: y = 16'h1ff;
			16'hc5a: y = 16'h1ff;
			16'hc5b: y = 16'h1ff;
			16'hc5c: y = 16'h1ff;
			16'hc5d: y = 16'h1ff;
			16'hc5e: y = 16'h1ff;
			16'hc5f: y = 16'h1ff;
			16'hc60: y = 16'h1ff;
			16'hc61: y = 16'h1ff;
			16'hc62: y = 16'h1ff;
			16'hc63: y = 16'h1ff;
			16'hc64: y = 16'h1ff;
			16'hc65: y = 16'h1ff;
			16'hc66: y = 16'h1ff;
			16'hc67: y = 16'h1ff;
			16'hc68: y = 16'h1ff;
			16'hc69: y = 16'h1ff;
			16'hc6a: y = 16'h1ff;
			16'hc6b: y = 16'h1ff;
			16'hc6c: y = 16'h1ff;
			16'hc6d: y = 16'h1ff;
			16'hc6e: y = 16'h1ff;
			16'hc6f: y = 16'h1ff;
			16'hc70: y = 16'h1ff;
			16'hc71: y = 16'h1ff;
			16'hc72: y = 16'h1ff;
			16'hc73: y = 16'h1ff;
			16'hc74: y = 16'h1ff;
			16'hc75: y = 16'h1ff;
			16'hc76: y = 16'h1ff;
			16'hc77: y = 16'h1ff;
			16'hc78: y = 16'h1ff;
			16'hc79: y = 16'h1ff;
			16'hc7a: y = 16'h1ff;
			16'hc7b: y = 16'h1ff;
			16'hc7c: y = 16'h1ff;
			16'hc7d: y = 16'h1ff;
			16'hc7e: y = 16'h1ff;
			16'hc7f: y = 16'h1ff;
			16'hc80: y = 16'h1ff;
			16'hc81: y = 16'h1ff;
			16'hc82: y = 16'h1ff;
			16'hc83: y = 16'h1ff;
			16'hc84: y = 16'h1ff;
			16'hc85: y = 16'h1ff;
			16'hc86: y = 16'h1ff;
			16'hc87: y = 16'h1ff;
			16'hc88: y = 16'h1ff;
			16'hc89: y = 16'h1ff;
			16'hc8a: y = 16'h1ff;
			16'hc8b: y = 16'h1ff;
			16'hc8c: y = 16'h1ff;
			16'hc8d: y = 16'h1ff;
			16'hc8e: y = 16'h1ff;
			16'hc8f: y = 16'h1ff;
			16'hc90: y = 16'h1ff;
			16'hc91: y = 16'h1ff;
			16'hc92: y = 16'h1ff;
			16'hc93: y = 16'h1ff;
			16'hc94: y = 16'h1ff;
			16'hc95: y = 16'h1ff;
			16'hc96: y = 16'h1ff;
			16'hc97: y = 16'h1ff;
			16'hc98: y = 16'h1ff;
			16'hc99: y = 16'h1ff;
			16'hc9a: y = 16'h1ff;
			16'hc9b: y = 16'h1ff;
			16'hc9c: y = 16'h1ff;
			16'hc9d: y = 16'h1ff;
			16'hc9e: y = 16'h1ff;
			16'hc9f: y = 16'h1ff;
			16'hca0: y = 16'h1ff;
			16'hca1: y = 16'h1ff;
			16'hca2: y = 16'h1ff;
			16'hca3: y = 16'h1ff;
			16'hca4: y = 16'h1ff;
			16'hca5: y = 16'h1ff;
			16'hca6: y = 16'h1ff;
			16'hca7: y = 16'h1ff;
			16'hca8: y = 16'h1ff;
			16'hca9: y = 16'h1ff;
			16'hcaa: y = 16'h1ff;
			16'hcab: y = 16'h1ff;
			16'hcac: y = 16'h1ff;
			16'hcad: y = 16'h1ff;
			16'hcae: y = 16'h1ff;
			16'hcaf: y = 16'h1ff;
			16'hcb0: y = 16'h1ff;
			16'hcb1: y = 16'h1ff;
			16'hcb2: y = 16'h1ff;
			16'hcb3: y = 16'h1ff;
			16'hcb4: y = 16'h1ff;
			16'hcb5: y = 16'h1ff;
			16'hcb6: y = 16'h1ff;
			16'hcb7: y = 16'h1ff;
			16'hcb8: y = 16'h1ff;
			16'hcb9: y = 16'h1ff;
			16'hcba: y = 16'h1ff;
			16'hcbb: y = 16'h1ff;
			16'hcbc: y = 16'h1ff;
			16'hcbd: y = 16'h1ff;
			16'hcbe: y = 16'h1ff;
			16'hcbf: y = 16'h1ff;
			16'hcc0: y = 16'h1ff;
			16'hcc1: y = 16'h1ff;
			16'hcc2: y = 16'h1ff;
			16'hcc3: y = 16'h1ff;
			16'hcc4: y = 16'h1ff;
			16'hcc5: y = 16'h1ff;
			16'hcc6: y = 16'h1ff;
			16'hcc7: y = 16'h1ff;
			16'hcc8: y = 16'h1ff;
			16'hcc9: y = 16'h1ff;
			16'hcca: y = 16'h1ff;
			16'hccb: y = 16'h1ff;
			16'hccc: y = 16'h1ff;
			16'hccd: y = 16'h1ff;
			16'hcce: y = 16'h1ff;
			16'hccf: y = 16'h1ff;
			16'hcd0: y = 16'h1ff;
			16'hcd1: y = 16'h1ff;
			16'hcd2: y = 16'h1ff;
			16'hcd3: y = 16'h1ff;
			16'hcd4: y = 16'h1ff;
			16'hcd5: y = 16'h1ff;
			16'hcd6: y = 16'h1ff;
			16'hcd7: y = 16'h1ff;
			16'hcd8: y = 16'h1ff;
			16'hcd9: y = 16'h1ff;
			16'hcda: y = 16'h1ff;
			16'hcdb: y = 16'h1ff;
			16'hcdc: y = 16'h1ff;
			16'hcdd: y = 16'h1ff;
			16'hcde: y = 16'h1ff;
			16'hcdf: y = 16'h1ff;
			16'hce0: y = 16'h1ff;
			16'hce1: y = 16'h1ff;
			16'hce2: y = 16'h1ff;
			16'hce3: y = 16'h1ff;
			16'hce4: y = 16'h1ff;
			16'hce5: y = 16'h1ff;
			16'hce6: y = 16'h1ff;
			16'hce7: y = 16'h1ff;
			16'hce8: y = 16'h1ff;
			16'hce9: y = 16'h1ff;
			16'hcea: y = 16'h1ff;
			16'hceb: y = 16'h1ff;
			16'hcec: y = 16'h1ff;
			16'hced: y = 16'h1ff;
			16'hcee: y = 16'h1ff;
			16'hcef: y = 16'h1ff;
			16'hcf0: y = 16'h1ff;
			16'hcf1: y = 16'h1ff;
			16'hcf2: y = 16'h1ff;
			16'hcf3: y = 16'h1ff;
			16'hcf4: y = 16'h1ff;
			16'hcf5: y = 16'h1ff;
			16'hcf6: y = 16'h1ff;
			16'hcf7: y = 16'h1ff;
			16'hcf8: y = 16'h1ff;
			16'hcf9: y = 16'h1ff;
			16'hcfa: y = 16'h1ff;
			16'hcfb: y = 16'h1ff;
			16'hcfc: y = 16'h1ff;
			16'hcfd: y = 16'h1ff;
			16'hcfe: y = 16'h1ff;
			16'hcff: y = 16'h1ff;
			16'hd00: y = 16'h1ff;
			16'hd01: y = 16'h1ff;
			16'hd02: y = 16'h1ff;
			16'hd03: y = 16'h1ff;
			16'hd04: y = 16'h1ff;
			16'hd05: y = 16'h1ff;
			16'hd06: y = 16'h1ff;
			16'hd07: y = 16'h1ff;
			16'hd08: y = 16'h1ff;
			16'hd09: y = 16'h1ff;
			16'hd0a: y = 16'h1ff;
			16'hd0b: y = 16'h1ff;
			16'hd0c: y = 16'h1ff;
			16'hd0d: y = 16'h1ff;
			16'hd0e: y = 16'h1ff;
			16'hd0f: y = 16'h1ff;
			16'hd10: y = 16'h1ff;
			16'hd11: y = 16'h1ff;
			16'hd12: y = 16'h1ff;
			16'hd13: y = 16'h1ff;
			16'hd14: y = 16'h1ff;
			16'hd15: y = 16'h1ff;
			16'hd16: y = 16'h1ff;
			16'hd17: y = 16'h1ff;
			16'hd18: y = 16'h1ff;
			16'hd19: y = 16'h1ff;
			16'hd1a: y = 16'h1ff;
			16'hd1b: y = 16'h1ff;
			16'hd1c: y = 16'h1ff;
			16'hd1d: y = 16'h1ff;
			16'hd1e: y = 16'h1ff;
			16'hd1f: y = 16'h1ff;
			16'hd20: y = 16'h1ff;
			16'hd21: y = 16'h1ff;
			16'hd22: y = 16'h1ff;
			16'hd23: y = 16'h1ff;
			16'hd24: y = 16'h1ff;
			16'hd25: y = 16'h1ff;
			16'hd26: y = 16'h1ff;
			16'hd27: y = 16'h1ff;
			16'hd28: y = 16'h1ff;
			16'hd29: y = 16'h1ff;
			16'hd2a: y = 16'h1ff;
			16'hd2b: y = 16'h1ff;
			16'hd2c: y = 16'h1ff;
			16'hd2d: y = 16'h1ff;
			16'hd2e: y = 16'h1ff;
			16'hd2f: y = 16'h1ff;
			16'hd30: y = 16'h1ff;
			16'hd31: y = 16'h1ff;
			16'hd32: y = 16'h1ff;
			16'hd33: y = 16'h1ff;
			16'hd34: y = 16'h1ff;
			16'hd35: y = 16'h1ff;
			16'hd36: y = 16'h1ff;
			16'hd37: y = 16'h1ff;
			16'hd38: y = 16'h1ff;
			16'hd39: y = 16'h1ff;
			16'hd3a: y = 16'h1ff;
			16'hd3b: y = 16'h1ff;
			16'hd3c: y = 16'h1ff;
			16'hd3d: y = 16'h1ff;
			16'hd3e: y = 16'h1ff;
			16'hd3f: y = 16'h1ff;
			16'hd40: y = 16'h1ff;
			16'hd41: y = 16'h1ff;
			16'hd42: y = 16'h1ff;
			16'hd43: y = 16'h1ff;
			16'hd44: y = 16'h1ff;
			16'hd45: y = 16'h1ff;
			16'hd46: y = 16'h1ff;
			16'hd47: y = 16'h1ff;
			16'hd48: y = 16'h1ff;
			16'hd49: y = 16'h1ff;
			16'hd4a: y = 16'h1ff;
			16'hd4b: y = 16'h1ff;
			16'hd4c: y = 16'h1ff;
			16'hd4d: y = 16'h1ff;
			16'hd4e: y = 16'h1ff;
			16'hd4f: y = 16'h1ff;
			16'hd50: y = 16'h1ff;
			16'hd51: y = 16'h1ff;
			16'hd52: y = 16'h1ff;
			16'hd53: y = 16'h1ff;
			16'hd54: y = 16'h1ff;
			16'hd55: y = 16'h1ff;
			16'hd56: y = 16'h1ff;
			16'hd57: y = 16'h1ff;
			16'hd58: y = 16'h1ff;
			16'hd59: y = 16'h1ff;
			16'hd5a: y = 16'h1ff;
			16'hd5b: y = 16'h1ff;
			16'hd5c: y = 16'h1ff;
			16'hd5d: y = 16'h1ff;
			16'hd5e: y = 16'h1ff;
			16'hd5f: y = 16'h1ff;
			16'hd60: y = 16'h1ff;
			16'hd61: y = 16'h1ff;
			16'hd62: y = 16'h1ff;
			16'hd63: y = 16'h1ff;
			16'hd64: y = 16'h1ff;
			16'hd65: y = 16'h1ff;
			16'hd66: y = 16'h1ff;
			16'hd67: y = 16'h1ff;
			16'hd68: y = 16'h1ff;
			16'hd69: y = 16'h1ff;
			16'hd6a: y = 16'h1ff;
			16'hd6b: y = 16'h1ff;
			16'hd6c: y = 16'h1ff;
			16'hd6d: y = 16'h1ff;
			16'hd6e: y = 16'h1ff;
			16'hd6f: y = 16'h1ff;
			16'hd70: y = 16'h1ff;
			16'hd71: y = 16'h1ff;
			16'hd72: y = 16'h1ff;
			16'hd73: y = 16'h1ff;
			16'hd74: y = 16'h1ff;
			16'hd75: y = 16'h1ff;
			16'hd76: y = 16'h1ff;
			16'hd77: y = 16'h1ff;
			16'hd78: y = 16'h1ff;
			16'hd79: y = 16'h1ff;
			16'hd7a: y = 16'h1ff;
			16'hd7b: y = 16'h1ff;
			16'hd7c: y = 16'h1ff;
			16'hd7d: y = 16'h1ff;
			16'hd7e: y = 16'h1ff;
			16'hd7f: y = 16'h1ff;
			16'hd80: y = 16'h1ff;
			16'hd81: y = 16'h1ff;
			16'hd82: y = 16'h1ff;
			16'hd83: y = 16'h1ff;
			16'hd84: y = 16'h1ff;
			16'hd85: y = 16'h1ff;
			16'hd86: y = 16'h1ff;
			16'hd87: y = 16'h1ff;
			16'hd88: y = 16'h1ff;
			16'hd89: y = 16'h1ff;
			16'hd8a: y = 16'h1ff;
			16'hd8b: y = 16'h1ff;
			16'hd8c: y = 16'h1ff;
			16'hd8d: y = 16'h1ff;
			16'hd8e: y = 16'h1ff;
			16'hd8f: y = 16'h1ff;
			16'hd90: y = 16'h1ff;
			16'hd91: y = 16'h1ff;
			16'hd92: y = 16'h1ff;
			16'hd93: y = 16'h1ff;
			16'hd94: y = 16'h1ff;
			16'hd95: y = 16'h1ff;
			16'hd96: y = 16'h1ff;
			16'hd97: y = 16'h1ff;
			16'hd98: y = 16'h1ff;
			16'hd99: y = 16'h1ff;
			16'hd9a: y = 16'h1ff;
			16'hd9b: y = 16'h1ff;
			16'hd9c: y = 16'h1ff;
			16'hd9d: y = 16'h1ff;
			16'hd9e: y = 16'h1ff;
			16'hd9f: y = 16'h1ff;
			16'hda0: y = 16'h1ff;
			16'hda1: y = 16'h1ff;
			16'hda2: y = 16'h1ff;
			16'hda3: y = 16'h1ff;
			16'hda4: y = 16'h1ff;
			16'hda5: y = 16'h1ff;
			16'hda6: y = 16'h1ff;
			16'hda7: y = 16'h1ff;
			16'hda8: y = 16'h1ff;
			16'hda9: y = 16'h1ff;
			16'hdaa: y = 16'h1ff;
			16'hdab: y = 16'h1ff;
			16'hdac: y = 16'h1ff;
			16'hdad: y = 16'h1ff;
			16'hdae: y = 16'h1ff;
			16'hdaf: y = 16'h1ff;
			16'hdb0: y = 16'h1ff;
			16'hdb1: y = 16'h1ff;
			16'hdb2: y = 16'h1ff;
			16'hdb3: y = 16'h1ff;
			16'hdb4: y = 16'h1ff;
			16'hdb5: y = 16'h1ff;
			16'hdb6: y = 16'h1ff;
			16'hdb7: y = 16'h1ff;
			16'hdb8: y = 16'h1ff;
			16'hdb9: y = 16'h1ff;
			16'hdba: y = 16'h1ff;
			16'hdbb: y = 16'h1ff;
			16'hdbc: y = 16'h1ff;
			16'hdbd: y = 16'h1ff;
			16'hdbe: y = 16'h1ff;
			16'hdbf: y = 16'h1ff;
			16'hdc0: y = 16'h1ff;
			16'hdc1: y = 16'h1ff;
			16'hdc2: y = 16'h1ff;
			16'hdc3: y = 16'h1ff;
			16'hdc4: y = 16'h1ff;
			16'hdc5: y = 16'h1ff;
			16'hdc6: y = 16'h1ff;
			16'hdc7: y = 16'h1ff;
			16'hdc8: y = 16'h1ff;
			16'hdc9: y = 16'h1ff;
			16'hdca: y = 16'h1ff;
			16'hdcb: y = 16'h1ff;
			16'hdcc: y = 16'h1ff;
			16'hdcd: y = 16'h1ff;
			16'hdce: y = 16'h1ff;
			16'hdcf: y = 16'h1ff;
			16'hdd0: y = 16'h1ff;
			16'hdd1: y = 16'h1ff;
			16'hdd2: y = 16'h1ff;
			16'hdd3: y = 16'h1ff;
			16'hdd4: y = 16'h1ff;
			16'hdd5: y = 16'h1ff;
			16'hdd6: y = 16'h1ff;
			16'hdd7: y = 16'h1ff;
			16'hdd8: y = 16'h1ff;
			16'hdd9: y = 16'h1ff;
			16'hdda: y = 16'h1ff;
			16'hddb: y = 16'h1ff;
			16'hddc: y = 16'h1ff;
			16'hddd: y = 16'h1ff;
			16'hdde: y = 16'h1ff;
			16'hddf: y = 16'h1ff;
			16'hde0: y = 16'h1ff;
			16'hde1: y = 16'h1ff;
			16'hde2: y = 16'h1ff;
			16'hde3: y = 16'h1ff;
			16'hde4: y = 16'h1ff;
			16'hde5: y = 16'h1ff;
			16'hde6: y = 16'h1ff;
			16'hde7: y = 16'h1ff;
			16'hde8: y = 16'h1ff;
			16'hde9: y = 16'h1ff;
			16'hdea: y = 16'h1ff;
			16'hdeb: y = 16'h1ff;
			16'hdec: y = 16'h1ff;
			16'hded: y = 16'h1ff;
			16'hdee: y = 16'h1ff;
			16'hdef: y = 16'h1ff;
			16'hdf0: y = 16'h1ff;
			16'hdf1: y = 16'h1ff;
			16'hdf2: y = 16'h1ff;
			16'hdf3: y = 16'h1ff;
			16'hdf4: y = 16'h1ff;
			16'hdf5: y = 16'h1ff;
			16'hdf6: y = 16'h1ff;
			16'hdf7: y = 16'h1ff;
			16'hdf8: y = 16'h1ff;
			16'hdf9: y = 16'h1ff;
			16'hdfa: y = 16'h1ff;
			16'hdfb: y = 16'h1ff;
			16'hdfc: y = 16'h1ff;
			16'hdfd: y = 16'h1ff;
			16'hdfe: y = 16'h1ff;
			16'hdff: y = 16'h1ff;
			16'he00: y = 16'h1ff;
			16'he01: y = 16'h1ff;
			16'he02: y = 16'h1ff;
			16'he03: y = 16'h1ff;
			16'he04: y = 16'h1ff;
			16'he05: y = 16'h1ff;
			16'he06: y = 16'h1ff;
			16'he07: y = 16'h1ff;
			16'he08: y = 16'h1ff;
			16'he09: y = 16'h1ff;
			16'he0a: y = 16'h1ff;
			16'he0b: y = 16'h1ff;
			16'he0c: y = 16'h1ff;
			16'he0d: y = 16'h1ff;
			16'he0e: y = 16'h1ff;
			16'he0f: y = 16'h1ff;
			16'he10: y = 16'h1ff;
			16'he11: y = 16'h1ff;
			16'he12: y = 16'h1ff;
			16'he13: y = 16'h1ff;
			16'he14: y = 16'h1ff;
			16'he15: y = 16'h1ff;
			16'he16: y = 16'h1ff;
			16'he17: y = 16'h1ff;
			16'he18: y = 16'h1ff;
			16'he19: y = 16'h1ff;
			16'he1a: y = 16'h1ff;
			16'he1b: y = 16'h1ff;
			16'he1c: y = 16'h1ff;
			16'he1d: y = 16'h1ff;
			16'he1e: y = 16'h1ff;
			16'he1f: y = 16'h1ff;
			16'he20: y = 16'h1ff;
			16'he21: y = 16'h1ff;
			16'he22: y = 16'h1ff;
			16'he23: y = 16'h1ff;
			16'he24: y = 16'h1ff;
			16'he25: y = 16'h1ff;
			16'he26: y = 16'h1ff;
			16'he27: y = 16'h1ff;
			16'he28: y = 16'h1ff;
			16'he29: y = 16'h1ff;
			16'he2a: y = 16'h1ff;
			16'he2b: y = 16'h1ff;
			16'he2c: y = 16'h1ff;
			16'he2d: y = 16'h1ff;
			16'he2e: y = 16'h1ff;
			16'he2f: y = 16'h1ff;
			16'he30: y = 16'h1ff;
			16'he31: y = 16'h1ff;
			16'he32: y = 16'h1ff;
			16'he33: y = 16'h1ff;
			16'he34: y = 16'h1ff;
			16'he35: y = 16'h1ff;
			16'he36: y = 16'h1ff;
			16'he37: y = 16'h1ff;
			16'he38: y = 16'h1ff;
			16'he39: y = 16'h1ff;
			16'he3a: y = 16'h1ff;
			16'he3b: y = 16'h1ff;
			16'he3c: y = 16'h1ff;
			16'he3d: y = 16'h1ff;
			16'he3e: y = 16'h1ff;
			16'he3f: y = 16'h1ff;
			16'he40: y = 16'h1ff;
			16'he41: y = 16'h1ff;
			16'he42: y = 16'h1ff;
			16'he43: y = 16'h1ff;
			16'he44: y = 16'h1ff;
			16'he45: y = 16'h1ff;
			16'he46: y = 16'h1ff;
			16'he47: y = 16'h1ff;
			16'he48: y = 16'h1ff;
			16'he49: y = 16'h1ff;
			16'he4a: y = 16'h1ff;
			16'he4b: y = 16'h1ff;
			16'he4c: y = 16'h1ff;
			16'he4d: y = 16'h1ff;
			16'he4e: y = 16'h1ff;
			16'he4f: y = 16'h1ff;
			16'he50: y = 16'h1ff;
			16'he51: y = 16'h1ff;
			16'he52: y = 16'h1ff;
			16'he53: y = 16'h1ff;
			16'he54: y = 16'h1ff;
			16'he55: y = 16'h1ff;
			16'he56: y = 16'h1ff;
			16'he57: y = 16'h1ff;
			16'he58: y = 16'h1ff;
			16'he59: y = 16'h1ff;
			16'he5a: y = 16'h1ff;
			16'he5b: y = 16'h1ff;
			16'he5c: y = 16'h1ff;
			16'he5d: y = 16'h1ff;
			16'he5e: y = 16'h1ff;
			16'he5f: y = 16'h1ff;
			16'he60: y = 16'h1ff;
			16'he61: y = 16'h1ff;
			16'he62: y = 16'h1ff;
			16'he63: y = 16'h1ff;
			16'he64: y = 16'h1ff;
			16'he65: y = 16'h1ff;
			16'he66: y = 16'h1ff;
			16'he67: y = 16'h1ff;
			16'he68: y = 16'h1ff;
			16'he69: y = 16'h1ff;
			16'he6a: y = 16'h1ff;
			16'he6b: y = 16'h1ff;
			16'he6c: y = 16'h1ff;
			16'he6d: y = 16'h1ff;
			16'he6e: y = 16'h1ff;
			16'he6f: y = 16'h1ff;
			16'he70: y = 16'h1ff;
			16'he71: y = 16'h1ff;
			16'he72: y = 16'h1ff;
			16'he73: y = 16'h1ff;
			16'he74: y = 16'h1ff;
			16'he75: y = 16'h1ff;
			16'he76: y = 16'h1ff;
			16'he77: y = 16'h1ff;
			16'he78: y = 16'h1ff;
			16'he79: y = 16'h1ff;
			16'he7a: y = 16'h1ff;
			16'he7b: y = 16'h1ff;
			16'he7c: y = 16'h1ff;
			16'he7d: y = 16'h1ff;
			16'he7e: y = 16'h1ff;
			16'he7f: y = 16'h1ff;
			16'he80: y = 16'h1ff;
			16'he81: y = 16'h1ff;
			16'he82: y = 16'h1ff;
			16'he83: y = 16'h1ff;
			16'he84: y = 16'h1ff;
			16'he85: y = 16'h1ff;
			16'he86: y = 16'h1ff;
			16'he87: y = 16'h1ff;
			16'he88: y = 16'h1ff;
			16'he89: y = 16'h1ff;
			16'he8a: y = 16'h1ff;
			16'he8b: y = 16'h1ff;
			16'he8c: y = 16'h1ff;
			16'he8d: y = 16'h1ff;
			16'he8e: y = 16'h1ff;
			16'he8f: y = 16'h1ff;
			16'he90: y = 16'h1ff;
			16'he91: y = 16'h1ff;
			16'he92: y = 16'h1ff;
			16'he93: y = 16'h1ff;
			16'he94: y = 16'h1ff;
			16'he95: y = 16'h1ff;
			16'he96: y = 16'h1ff;
			16'he97: y = 16'h1ff;
			16'he98: y = 16'h1ff;
			16'he99: y = 16'h1ff;
			16'he9a: y = 16'h1ff;
			16'he9b: y = 16'h1ff;
			16'he9c: y = 16'h1ff;
			16'he9d: y = 16'h1ff;
			16'he9e: y = 16'h1ff;
			16'he9f: y = 16'h1ff;
			16'hea0: y = 16'h1ff;
			16'hea1: y = 16'h1ff;
			16'hea2: y = 16'h1ff;
			16'hea3: y = 16'h1ff;
			16'hea4: y = 16'h1ff;
			16'hea5: y = 16'h1ff;
			16'hea6: y = 16'h1ff;
			16'hea7: y = 16'h1ff;
			16'hea8: y = 16'h1ff;
			16'hea9: y = 16'h1ff;
			16'heaa: y = 16'h1ff;
			16'heab: y = 16'h1ff;
			16'heac: y = 16'h1ff;
			16'head: y = 16'h1ff;
			16'heae: y = 16'h1ff;
			16'heaf: y = 16'h1ff;
			16'heb0: y = 16'h1ff;
			16'heb1: y = 16'h1ff;
			16'heb2: y = 16'h1ff;
			16'heb3: y = 16'h1ff;
			16'heb4: y = 16'h1ff;
			16'heb5: y = 16'h1ff;
			16'heb6: y = 16'h1ff;
			16'heb7: y = 16'h1ff;
			16'heb8: y = 16'h1ff;
			16'heb9: y = 16'h1ff;
			16'heba: y = 16'h1ff;
			16'hebb: y = 16'h1ff;
			16'hebc: y = 16'h1ff;
			16'hebd: y = 16'h1ff;
			16'hebe: y = 16'h1ff;
			16'hebf: y = 16'h1ff;
			16'hec0: y = 16'h1ff;
			16'hec1: y = 16'h1ff;
			16'hec2: y = 16'h1ff;
			16'hec3: y = 16'h1ff;
			16'hec4: y = 16'h1ff;
			16'hec5: y = 16'h1ff;
			16'hec6: y = 16'h1ff;
			16'hec7: y = 16'h1ff;
			16'hec8: y = 16'h1ff;
			16'hec9: y = 16'h1ff;
			16'heca: y = 16'h1ff;
			16'hecb: y = 16'h1ff;
			16'hecc: y = 16'h1ff;
			16'hecd: y = 16'h1ff;
			16'hece: y = 16'h1ff;
			16'hecf: y = 16'h1ff;
			16'hed0: y = 16'h1ff;
			16'hed1: y = 16'h1ff;
			16'hed2: y = 16'h1ff;
			16'hed3: y = 16'h1ff;
			16'hed4: y = 16'h1ff;
			16'hed5: y = 16'h1ff;
			16'hed6: y = 16'h1ff;
			16'hed7: y = 16'h1ff;
			16'hed8: y = 16'h1ff;
			16'hed9: y = 16'h1ff;
			16'heda: y = 16'h1ff;
			16'hedb: y = 16'h1ff;
			16'hedc: y = 16'h1ff;
			16'hedd: y = 16'h1ff;
			16'hede: y = 16'h1ff;
			16'hedf: y = 16'h1ff;
			16'hee0: y = 16'h1ff;
			16'hee1: y = 16'h1ff;
			16'hee2: y = 16'h1ff;
			16'hee3: y = 16'h1ff;
			16'hee4: y = 16'h1ff;
			16'hee5: y = 16'h1ff;
			16'hee6: y = 16'h1ff;
			16'hee7: y = 16'h1ff;
			16'hee8: y = 16'h1ff;
			16'hee9: y = 16'h1ff;
			16'heea: y = 16'h1ff;
			16'heeb: y = 16'h1ff;
			16'heec: y = 16'h1ff;
			16'heed: y = 16'h1ff;
			16'heee: y = 16'h1ff;
			16'heef: y = 16'h1ff;
			16'hef0: y = 16'h1ff;
			16'hef1: y = 16'h1ff;
			16'hef2: y = 16'h1ff;
			16'hef3: y = 16'h1ff;
			16'hef4: y = 16'h1ff;
			16'hef5: y = 16'h1ff;
			16'hef6: y = 16'h1ff;
			16'hef7: y = 16'h1ff;
			16'hef8: y = 16'h1ff;
			16'hef9: y = 16'h1ff;
			16'hefa: y = 16'h1ff;
			16'hefb: y = 16'h1ff;
			16'hefc: y = 16'h1ff;
			16'hefd: y = 16'h1ff;
			16'hefe: y = 16'h1ff;
			16'heff: y = 16'h1ff;
			16'hf00: y = 16'h1ff;
			16'hf01: y = 16'h1ff;
			16'hf02: y = 16'h1ff;
			16'hf03: y = 16'h1ff;
			16'hf04: y = 16'h1ff;
			16'hf05: y = 16'h1ff;
			16'hf06: y = 16'h1ff;
			16'hf07: y = 16'h1ff;
			16'hf08: y = 16'h1ff;
			16'hf09: y = 16'h1ff;
			16'hf0a: y = 16'h1ff;
			16'hf0b: y = 16'h1ff;
			16'hf0c: y = 16'h1ff;
			16'hf0d: y = 16'h1ff;
			16'hf0e: y = 16'h1ff;
			16'hf0f: y = 16'h1ff;
			16'hf10: y = 16'h1ff;
			16'hf11: y = 16'h1ff;
			16'hf12: y = 16'h1ff;
			16'hf13: y = 16'h1ff;
			16'hf14: y = 16'h1ff;
			16'hf15: y = 16'h1ff;
			16'hf16: y = 16'h1ff;
			16'hf17: y = 16'h1ff;
			16'hf18: y = 16'h1ff;
			16'hf19: y = 16'h1ff;
			16'hf1a: y = 16'h1ff;
			16'hf1b: y = 16'h1ff;
			16'hf1c: y = 16'h1ff;
			16'hf1d: y = 16'h1ff;
			16'hf1e: y = 16'h1ff;
			16'hf1f: y = 16'h1ff;
			16'hf20: y = 16'h1ff;
			16'hf21: y = 16'h1ff;
			16'hf22: y = 16'h1ff;
			16'hf23: y = 16'h1ff;
			16'hf24: y = 16'h1ff;
			16'hf25: y = 16'h1ff;
			16'hf26: y = 16'h1ff;
			16'hf27: y = 16'h1ff;
			16'hf28: y = 16'h1ff;
			16'hf29: y = 16'h1ff;
			16'hf2a: y = 16'h1ff;
			16'hf2b: y = 16'h1ff;
			16'hf2c: y = 16'h1ff;
			16'hf2d: y = 16'h1ff;
			16'hf2e: y = 16'h1ff;
			16'hf2f: y = 16'h1ff;
			16'hf30: y = 16'h1ff;
			16'hf31: y = 16'h1ff;
			16'hf32: y = 16'h1ff;
			16'hf33: y = 16'h1ff;
			16'hf34: y = 16'h1ff;
			16'hf35: y = 16'h1ff;
			16'hf36: y = 16'h1ff;
			16'hf37: y = 16'h1ff;
			16'hf38: y = 16'h1ff;
			16'hf39: y = 16'h1ff;
			16'hf3a: y = 16'h1ff;
			16'hf3b: y = 16'h1ff;
			16'hf3c: y = 16'h1ff;
			16'hf3d: y = 16'h1ff;
			16'hf3e: y = 16'h1ff;
			16'hf3f: y = 16'h1ff;
			16'hf40: y = 16'h1ff;
			16'hf41: y = 16'h1ff;
			16'hf42: y = 16'h1ff;
			16'hf43: y = 16'h1ff;
			16'hf44: y = 16'h1ff;
			16'hf45: y = 16'h1ff;
			16'hf46: y = 16'h1ff;
			16'hf47: y = 16'h1ff;
			16'hf48: y = 16'h1ff;
			16'hf49: y = 16'h1ff;
			16'hf4a: y = 16'h1ff;
			16'hf4b: y = 16'h1ff;
			16'hf4c: y = 16'h1ff;
			16'hf4d: y = 16'h1ff;
			16'hf4e: y = 16'h1ff;
			16'hf4f: y = 16'h1ff;
			16'hf50: y = 16'h1ff;
			16'hf51: y = 16'h1ff;
			16'hf52: y = 16'h1ff;
			16'hf53: y = 16'h1ff;
			16'hf54: y = 16'h1ff;
			16'hf55: y = 16'h1ff;
			16'hf56: y = 16'h1ff;
			16'hf57: y = 16'h1ff;
			16'hf58: y = 16'h1ff;
			16'hf59: y = 16'h1ff;
			16'hf5a: y = 16'h1ff;
			16'hf5b: y = 16'h1ff;
			16'hf5c: y = 16'h1ff;
			16'hf5d: y = 16'h1ff;
			16'hf5e: y = 16'h1ff;
			16'hf5f: y = 16'h1ff;
			16'hf60: y = 16'h1ff;
			16'hf61: y = 16'h1ff;
			16'hf62: y = 16'h1ff;
			16'hf63: y = 16'h1ff;
			16'hf64: y = 16'h1ff;
			16'hf65: y = 16'h1ff;
			16'hf66: y = 16'h1ff;
			16'hf67: y = 16'h1ff;
			16'hf68: y = 16'h1ff;
			16'hf69: y = 16'h1ff;
			16'hf6a: y = 16'h1ff;
			16'hf6b: y = 16'h1ff;
			16'hf6c: y = 16'h1ff;
			16'hf6d: y = 16'h1ff;
			16'hf6e: y = 16'h1ff;
			16'hf6f: y = 16'h1ff;
			16'hf70: y = 16'h1ff;
			16'hf71: y = 16'h1ff;
			16'hf72: y = 16'h1ff;
			16'hf73: y = 16'h1ff;
			16'hf74: y = 16'h1ff;
			16'hf75: y = 16'h1ff;
			16'hf76: y = 16'h1ff;
			16'hf77: y = 16'h1ff;
			16'hf78: y = 16'h1ff;
			16'hf79: y = 16'h1ff;
			16'hf7a: y = 16'h1ff;
			16'hf7b: y = 16'h1ff;
			16'hf7c: y = 16'h1ff;
			16'hf7d: y = 16'h1ff;
			16'hf7e: y = 16'h1ff;
			16'hf7f: y = 16'h1ff;
			16'hf80: y = 16'h1ff;
			16'hf81: y = 16'h1ff;
			16'hf82: y = 16'h1ff;
			16'hf83: y = 16'h1ff;
			16'hf84: y = 16'h1ff;
			16'hf85: y = 16'h1ff;
			16'hf86: y = 16'h1ff;
			16'hf87: y = 16'h1ff;
			16'hf88: y = 16'h1ff;
			16'hf89: y = 16'h1ff;
			16'hf8a: y = 16'h1ff;
			16'hf8b: y = 16'h1ff;
			16'hf8c: y = 16'h1ff;
			16'hf8d: y = 16'h1ff;
			16'hf8e: y = 16'h1ff;
			16'hf8f: y = 16'h1ff;
			16'hf90: y = 16'h1ff;
			16'hf91: y = 16'h1ff;
			16'hf92: y = 16'h1ff;
			16'hf93: y = 16'h1ff;
			16'hf94: y = 16'h1ff;
			16'hf95: y = 16'h1ff;
			16'hf96: y = 16'h1ff;
			16'hf97: y = 16'h1ff;
			16'hf98: y = 16'h1ff;
			16'hf99: y = 16'h1ff;
			16'hf9a: y = 16'h1ff;
			16'hf9b: y = 16'h1ff;
			16'hf9c: y = 16'h1ff;
			16'hf9d: y = 16'h1ff;
			16'hf9e: y = 16'h1ff;
			16'hf9f: y = 16'h1ff;
			16'hfa0: y = 16'h1ff;
			16'hfa1: y = 16'h1ff;
			16'hfa2: y = 16'h1ff;
			16'hfa3: y = 16'h1ff;
			16'hfa4: y = 16'h1ff;
			16'hfa5: y = 16'h1ff;
			16'hfa6: y = 16'h1ff;
			16'hfa7: y = 16'h1ff;
			16'hfa8: y = 16'h1ff;
			16'hfa9: y = 16'h1ff;
			16'hfaa: y = 16'h1ff;
			16'hfab: y = 16'h1ff;
			16'hfac: y = 16'h1ff;
			16'hfad: y = 16'h1ff;
			16'hfae: y = 16'h1ff;
			16'hfaf: y = 16'h1ff;
			16'hfb0: y = 16'h1ff;
			16'hfb1: y = 16'h1ff;
			16'hfb2: y = 16'h1ff;
			16'hfb3: y = 16'h1ff;
			16'hfb4: y = 16'h1ff;
			16'hfb5: y = 16'h1ff;
			16'hfb6: y = 16'h1ff;
			16'hfb7: y = 16'h1ff;
			16'hfb8: y = 16'h1ff;
			16'hfb9: y = 16'h1ff;
			16'hfba: y = 16'h1ff;
			16'hfbb: y = 16'h1ff;
			16'hfbc: y = 16'h1ff;
			16'hfbd: y = 16'h1ff;
			16'hfbe: y = 16'h1ff;
			16'hfbf: y = 16'h1ff;
			16'hfc0: y = 16'h1ff;
			16'hfc1: y = 16'h1ff;
			16'hfc2: y = 16'h1ff;
			16'hfc3: y = 16'h1ff;
			16'hfc4: y = 16'h1ff;
			16'hfc5: y = 16'h1ff;
			16'hfc6: y = 16'h1ff;
			16'hfc7: y = 16'h1ff;
			16'hfc8: y = 16'h1ff;
			16'hfc9: y = 16'h1ff;
			16'hfca: y = 16'h1ff;
			16'hfcb: y = 16'h1ff;
			16'hfcc: y = 16'h1ff;
			16'hfcd: y = 16'h1ff;
			16'hfce: y = 16'h1ff;
			16'hfcf: y = 16'h1ff;
			16'hfd0: y = 16'h1ff;
			16'hfd1: y = 16'h1ff;
			16'hfd2: y = 16'h1ff;
			16'hfd3: y = 16'h1ff;
			16'hfd4: y = 16'h1ff;
			16'hfd5: y = 16'h1ff;
			16'hfd6: y = 16'h1ff;
			16'hfd7: y = 16'h1ff;
			16'hfd8: y = 16'h1ff;
			16'hfd9: y = 16'h1ff;
			16'hfda: y = 16'h1ff;
			16'hfdb: y = 16'h1ff;
			16'hfdc: y = 16'h1ff;
			16'hfdd: y = 16'h1ff;
			16'hfde: y = 16'h1ff;
			16'hfdf: y = 16'h1ff;
			16'hfe0: y = 16'h1ff;
			16'hfe1: y = 16'h1ff;
			16'hfe2: y = 16'h1ff;
			16'hfe3: y = 16'h1ff;
			16'hfe4: y = 16'h1ff;
			16'hfe5: y = 16'h1ff;
			16'hfe6: y = 16'h1ff;
			16'hfe7: y = 16'h1ff;
			16'hfe8: y = 16'h1ff;
			16'hfe9: y = 16'h1ff;
			16'hfea: y = 16'h1ff;
			16'hfeb: y = 16'h1ff;
			16'hfec: y = 16'h1ff;
			16'hfed: y = 16'h1ff;
			16'hfee: y = 16'h1ff;
			16'hfef: y = 16'h1ff;
			16'hff0: y = 16'h1ff;
			16'hff1: y = 16'h1ff;
			16'hff2: y = 16'h1ff;
			16'hff3: y = 16'h1ff;
			16'hff4: y = 16'h1ff;
			16'hff5: y = 16'h1ff;
			16'hff6: y = 16'h1ff;
			16'hff7: y = 16'h1ff;
			16'hff8: y = 16'h1ff;
			16'hff9: y = 16'h1ff;
			16'hffa: y = 16'h1ff;
			16'hffb: y = 16'h1ff;
			16'hffc: y = 16'h1ff;
			16'hffd: y = 16'h1ff;
			16'hffe: y = 16'h1ff;
			16'hfff: y = 16'h1ff;
			16'h1000: y = 16'h1ff;
			16'h1001: y = 16'h1ff;
			16'h1002: y = 16'h1ff;
			16'h1003: y = 16'h1ff;
			16'h1004: y = 16'h1ff;
			16'h1005: y = 16'h1ff;
			16'h1006: y = 16'h1ff;
			16'h1007: y = 16'h1ff;
			16'h1008: y = 16'h1ff;
			16'h1009: y = 16'h1ff;
			16'h100a: y = 16'h1ff;
			16'h100b: y = 16'h1ff;
			16'h100c: y = 16'h1ff;
			16'h100d: y = 16'h1ff;
			16'h100e: y = 16'h1ff;
			16'h100f: y = 16'h1ff;
			16'h1010: y = 16'h1ff;
			16'h1011: y = 16'h1ff;
			16'h1012: y = 16'h1ff;
			16'h1013: y = 16'h1ff;
			16'h1014: y = 16'h1ff;
			16'h1015: y = 16'h1ff;
			16'h1016: y = 16'h1ff;
			16'h1017: y = 16'h1ff;
			16'h1018: y = 16'h1ff;
			16'h1019: y = 16'h1ff;
			16'h101a: y = 16'h1ff;
			16'h101b: y = 16'h1ff;
			16'h101c: y = 16'h1ff;
			16'h101d: y = 16'h1ff;
			16'h101e: y = 16'h1ff;
			16'h101f: y = 16'h1ff;
			16'h1020: y = 16'h1ff;
			16'h1021: y = 16'h1ff;
			16'h1022: y = 16'h1ff;
			16'h1023: y = 16'h1ff;
			16'h1024: y = 16'h1ff;
			16'h1025: y = 16'h1ff;
			16'h1026: y = 16'h1ff;
			16'h1027: y = 16'h1ff;
			16'h1028: y = 16'h1ff;
			16'h1029: y = 16'h1ff;
			16'h102a: y = 16'h1ff;
			16'h102b: y = 16'h1ff;
			16'h102c: y = 16'h1ff;
			16'h102d: y = 16'h1ff;
			16'h102e: y = 16'h1ff;
			16'h102f: y = 16'h1ff;
			16'h1030: y = 16'h1ff;
			16'h1031: y = 16'h1ff;
			16'h1032: y = 16'h1ff;
			16'h1033: y = 16'h1ff;
			16'h1034: y = 16'h1ff;
			16'h1035: y = 16'h1ff;
			16'h1036: y = 16'h1ff;
			16'h1037: y = 16'h1ff;
			16'h1038: y = 16'h1ff;
			16'h1039: y = 16'h1ff;
			16'h103a: y = 16'h1ff;
			16'h103b: y = 16'h1ff;
			16'h103c: y = 16'h1ff;
			16'h103d: y = 16'h1ff;
			16'h103e: y = 16'h1ff;
			16'h103f: y = 16'h1ff;
			16'h1040: y = 16'h1ff;
			16'h1041: y = 16'h1ff;
			16'h1042: y = 16'h1ff;
			16'h1043: y = 16'h1ff;
			16'h1044: y = 16'h1ff;
			16'h1045: y = 16'h1ff;
			16'h1046: y = 16'h1ff;
			16'h1047: y = 16'h1ff;
			16'h1048: y = 16'h1ff;
			16'h1049: y = 16'h1ff;
			16'h104a: y = 16'h1ff;
			16'h104b: y = 16'h1ff;
			16'h104c: y = 16'h1ff;
			16'h104d: y = 16'h1ff;
			16'h104e: y = 16'h1ff;
			16'h104f: y = 16'h1ff;
			16'h1050: y = 16'h1ff;
			16'h1051: y = 16'h1ff;
			16'h1052: y = 16'h1ff;
			16'h1053: y = 16'h1ff;
			16'h1054: y = 16'h1ff;
			16'h1055: y = 16'h1ff;
			16'h1056: y = 16'h1ff;
			16'h1057: y = 16'h1ff;
			16'h1058: y = 16'h1ff;
			16'h1059: y = 16'h1ff;
			16'h105a: y = 16'h1ff;
			16'h105b: y = 16'h1ff;
			16'h105c: y = 16'h1ff;
			16'h105d: y = 16'h1ff;
			16'h105e: y = 16'h1ff;
			16'h105f: y = 16'h1ff;
			16'h1060: y = 16'h1ff;
			16'h1061: y = 16'h1ff;
			16'h1062: y = 16'h1ff;
			16'h1063: y = 16'h1ff;
			16'h1064: y = 16'h1ff;
			16'h1065: y = 16'h1ff;
			16'h1066: y = 16'h1ff;
			16'h1067: y = 16'h1ff;
			16'h1068: y = 16'h1ff;
			16'h1069: y = 16'h1ff;
			16'h106a: y = 16'h1ff;
			16'h106b: y = 16'h1ff;
			16'h106c: y = 16'h1ff;
			16'h106d: y = 16'h1ff;
			16'h106e: y = 16'h1ff;
			16'h106f: y = 16'h1ff;
			16'h1070: y = 16'h1ff;
			16'h1071: y = 16'h1ff;
			16'h1072: y = 16'h1ff;
			16'h1073: y = 16'h1ff;
			16'h1074: y = 16'h1ff;
			16'h1075: y = 16'h1ff;
			16'h1076: y = 16'h1ff;
			16'h1077: y = 16'h1ff;
			16'h1078: y = 16'h1ff;
			16'h1079: y = 16'h1ff;
			16'h107a: y = 16'h1ff;
			16'h107b: y = 16'h1ff;
			16'h107c: y = 16'h1ff;
			16'h107d: y = 16'h1ff;
			16'h107e: y = 16'h1ff;
			16'h107f: y = 16'h1ff;
			16'h1080: y = 16'h1ff;
			16'h1081: y = 16'h1ff;
			16'h1082: y = 16'h1ff;
			16'h1083: y = 16'h1ff;
			16'h1084: y = 16'h1ff;
			16'h1085: y = 16'h1ff;
			16'h1086: y = 16'h1ff;
			16'h1087: y = 16'h1ff;
			16'h1088: y = 16'h1ff;
			16'h1089: y = 16'h1ff;
			16'h108a: y = 16'h1ff;
			16'h108b: y = 16'h1ff;
			16'h108c: y = 16'h1ff;
			16'h108d: y = 16'h1ff;
			16'h108e: y = 16'h1ff;
			16'h108f: y = 16'h1ff;
			16'h1090: y = 16'h1ff;
			16'h1091: y = 16'h1ff;
			16'h1092: y = 16'h1ff;
			16'h1093: y = 16'h1ff;
			16'h1094: y = 16'h1ff;
			16'h1095: y = 16'h1ff;
			16'h1096: y = 16'h1ff;
			16'h1097: y = 16'h1ff;
			16'h1098: y = 16'h1ff;
			16'h1099: y = 16'h1ff;
			16'h109a: y = 16'h1ff;
			16'h109b: y = 16'h1ff;
			16'h109c: y = 16'h1ff;
			16'h109d: y = 16'h1ff;
			16'h109e: y = 16'h1ff;
			16'h109f: y = 16'h1ff;
			16'h10a0: y = 16'h1ff;
			16'h10a1: y = 16'h1ff;
			16'h10a2: y = 16'h1ff;
			16'h10a3: y = 16'h1ff;
			16'h10a4: y = 16'h1ff;
			16'h10a5: y = 16'h1ff;
			16'h10a6: y = 16'h1ff;
			16'h10a7: y = 16'h1ff;
			16'h10a8: y = 16'h1ff;
			16'h10a9: y = 16'h1ff;
			16'h10aa: y = 16'h1ff;
			16'h10ab: y = 16'h1ff;
			16'h10ac: y = 16'h1ff;
			16'h10ad: y = 16'h1ff;
			16'h10ae: y = 16'h1ff;
			16'h10af: y = 16'h1ff;
			16'h10b0: y = 16'h1ff;
			16'h10b1: y = 16'h1ff;
			16'h10b2: y = 16'h1ff;
			16'h10b3: y = 16'h1ff;
			16'h10b4: y = 16'h1ff;
			16'h10b5: y = 16'h1ff;
			16'h10b6: y = 16'h1ff;
			16'h10b7: y = 16'h1ff;
			16'h10b8: y = 16'h1ff;
			16'h10b9: y = 16'h1ff;
			16'h10ba: y = 16'h1ff;
			16'h10bb: y = 16'h1ff;
			16'h10bc: y = 16'h1ff;
			16'h10bd: y = 16'h1ff;
			16'h10be: y = 16'h1ff;
			16'h10bf: y = 16'h1ff;
			16'h10c0: y = 16'h1ff;
			16'h10c1: y = 16'h1ff;
			16'h10c2: y = 16'h1ff;
			16'h10c3: y = 16'h1ff;
			16'h10c4: y = 16'h1ff;
			16'h10c5: y = 16'h1ff;
			16'h10c6: y = 16'h1ff;
			16'h10c7: y = 16'h1ff;
			16'h10c8: y = 16'h1ff;
			16'h10c9: y = 16'h1ff;
			16'h10ca: y = 16'h1ff;
			16'h10cb: y = 16'h1ff;
			16'h10cc: y = 16'h1ff;
			16'h10cd: y = 16'h1ff;
			16'h10ce: y = 16'h1ff;
			16'h10cf: y = 16'h1ff;
			16'h10d0: y = 16'h1ff;
			16'h10d1: y = 16'h1ff;
			16'h10d2: y = 16'h1ff;
			16'h10d3: y = 16'h1ff;
			16'h10d4: y = 16'h1ff;
			16'h10d5: y = 16'h1ff;
			16'h10d6: y = 16'h1ff;
			16'h10d7: y = 16'h1ff;
			16'h10d8: y = 16'h1ff;
			16'h10d9: y = 16'h1ff;
			16'h10da: y = 16'h1ff;
			16'h10db: y = 16'h1ff;
			16'h10dc: y = 16'h1ff;
			16'h10dd: y = 16'h1ff;
			16'h10de: y = 16'h1ff;
			16'h10df: y = 16'h1ff;
			16'h10e0: y = 16'h1ff;
			16'h10e1: y = 16'h1ff;
			16'h10e2: y = 16'h1ff;
			16'h10e3: y = 16'h1ff;
			16'h10e4: y = 16'h1ff;
			16'h10e5: y = 16'h1ff;
			16'h10e6: y = 16'h1ff;
			16'h10e7: y = 16'h1ff;
			16'h10e8: y = 16'h1ff;
			16'h10e9: y = 16'h1ff;
			16'h10ea: y = 16'h1ff;
			16'h10eb: y = 16'h1ff;
			16'h10ec: y = 16'h1ff;
			16'h10ed: y = 16'h1ff;
			16'h10ee: y = 16'h1ff;
			16'h10ef: y = 16'h1ff;
			16'h10f0: y = 16'h1ff;
			16'h10f1: y = 16'h1ff;
			16'h10f2: y = 16'h1ff;
			16'h10f3: y = 16'h1ff;
			16'h10f4: y = 16'h1ff;
			16'h10f5: y = 16'h1ff;
			16'h10f6: y = 16'h1ff;
			16'h10f7: y = 16'h1ff;
			16'h10f8: y = 16'h1ff;
			16'h10f9: y = 16'h1ff;
			16'h10fa: y = 16'h1ff;
			16'h10fb: y = 16'h1ff;
			16'h10fc: y = 16'h1ff;
			16'h10fd: y = 16'h1ff;
			16'h10fe: y = 16'h1ff;
			16'h10ff: y = 16'h1ff;
			16'h1100: y = 16'h1ff;
			16'h1101: y = 16'h1ff;
			16'h1102: y = 16'h1ff;
			16'h1103: y = 16'h1ff;
			16'h1104: y = 16'h1ff;
			16'h1105: y = 16'h1ff;
			16'h1106: y = 16'h1ff;
			16'h1107: y = 16'h1ff;
			16'h1108: y = 16'h1ff;
			16'h1109: y = 16'h1ff;
			16'h110a: y = 16'h1ff;
			16'h110b: y = 16'h1ff;
			16'h110c: y = 16'h1ff;
			16'h110d: y = 16'h1ff;
			16'h110e: y = 16'h1ff;
			16'h110f: y = 16'h1ff;
			16'h1110: y = 16'h1ff;
			16'h1111: y = 16'h1ff;
			16'h1112: y = 16'h1ff;
			16'h1113: y = 16'h1ff;
			16'h1114: y = 16'h1ff;
			16'h1115: y = 16'h1ff;
			16'h1116: y = 16'h1ff;
			16'h1117: y = 16'h1ff;
			16'h1118: y = 16'h1ff;
			16'h1119: y = 16'h1ff;
			16'h111a: y = 16'h1ff;
			16'h111b: y = 16'h1ff;
			16'h111c: y = 16'h1ff;
			16'h111d: y = 16'h1ff;
			16'h111e: y = 16'h1ff;
			16'h111f: y = 16'h1ff;
			16'h1120: y = 16'h1ff;
			16'h1121: y = 16'h1ff;
			16'h1122: y = 16'h1ff;
			16'h1123: y = 16'h1ff;
			16'h1124: y = 16'h1ff;
			16'h1125: y = 16'h1ff;
			16'h1126: y = 16'h1ff;
			16'h1127: y = 16'h1ff;
			16'h1128: y = 16'h1ff;
			16'h1129: y = 16'h1ff;
			16'h112a: y = 16'h1ff;
			16'h112b: y = 16'h1ff;
			16'h112c: y = 16'h1ff;
			16'h112d: y = 16'h1ff;
			16'h112e: y = 16'h1ff;
			16'h112f: y = 16'h1ff;
			16'h1130: y = 16'h1ff;
			16'h1131: y = 16'h1ff;
			16'h1132: y = 16'h1ff;
			16'h1133: y = 16'h1ff;
			16'h1134: y = 16'h1ff;
			16'h1135: y = 16'h1ff;
			16'h1136: y = 16'h1ff;
			16'h1137: y = 16'h1ff;
			16'h1138: y = 16'h1ff;
			16'h1139: y = 16'h1ff;
			16'h113a: y = 16'h1ff;
			16'h113b: y = 16'h1ff;
			16'h113c: y = 16'h1ff;
			16'h113d: y = 16'h1ff;
			16'h113e: y = 16'h1ff;
			16'h113f: y = 16'h1ff;
			16'h1140: y = 16'h1ff;
			16'h1141: y = 16'h1ff;
			16'h1142: y = 16'h1ff;
			16'h1143: y = 16'h1ff;
			16'h1144: y = 16'h1ff;
			16'h1145: y = 16'h1ff;
			16'h1146: y = 16'h1ff;
			16'h1147: y = 16'h1ff;
			16'h1148: y = 16'h1ff;
			16'h1149: y = 16'h1ff;
			16'h114a: y = 16'h1ff;
			16'h114b: y = 16'h1ff;
			16'h114c: y = 16'h1ff;
			16'h114d: y = 16'h1ff;
			16'h114e: y = 16'h1ff;
			16'h114f: y = 16'h1ff;
			16'h1150: y = 16'h1ff;
			16'h1151: y = 16'h1ff;
			16'h1152: y = 16'h1ff;
			16'h1153: y = 16'h1ff;
			16'h1154: y = 16'h1ff;
			16'h1155: y = 16'h1ff;
			16'h1156: y = 16'h1ff;
			16'h1157: y = 16'h1ff;
			16'h1158: y = 16'h1ff;
			16'h1159: y = 16'h1ff;
			16'h115a: y = 16'h1ff;
			16'h115b: y = 16'h1ff;
			16'h115c: y = 16'h1ff;
			16'h115d: y = 16'h1ff;
			16'h115e: y = 16'h1ff;
			16'h115f: y = 16'h1ff;
			16'h1160: y = 16'h1ff;
			16'h1161: y = 16'h1ff;
			16'h1162: y = 16'h1ff;
			16'h1163: y = 16'h1ff;
			16'h1164: y = 16'h1ff;
			16'h1165: y = 16'h1ff;
			16'h1166: y = 16'h1ff;
			16'h1167: y = 16'h1ff;
			16'h1168: y = 16'h1ff;
			16'h1169: y = 16'h1ff;
			16'h116a: y = 16'h1ff;
			16'h116b: y = 16'h1ff;
			16'h116c: y = 16'h1ff;
			16'h116d: y = 16'h1ff;
			16'h116e: y = 16'h1ff;
			16'h116f: y = 16'h1ff;
			16'h1170: y = 16'h1ff;
			16'h1171: y = 16'h1ff;
			16'h1172: y = 16'h1ff;
			16'h1173: y = 16'h1ff;
			16'h1174: y = 16'h1ff;
			16'h1175: y = 16'h1ff;
			16'h1176: y = 16'h1ff;
			16'h1177: y = 16'h1ff;
			16'h1178: y = 16'h1ff;
			16'h1179: y = 16'h1ff;
			16'h117a: y = 16'h1ff;
			16'h117b: y = 16'h1ff;
			16'h117c: y = 16'h1ff;
			16'h117d: y = 16'h1ff;
			16'h117e: y = 16'h1ff;
			16'h117f: y = 16'h1ff;
			16'h1180: y = 16'h1ff;
			16'h1181: y = 16'h1ff;
			16'h1182: y = 16'h1ff;
			16'h1183: y = 16'h1ff;
			16'h1184: y = 16'h1ff;
			16'h1185: y = 16'h1ff;
			16'h1186: y = 16'h1ff;
			16'h1187: y = 16'h1ff;
			16'h1188: y = 16'h1ff;
			16'h1189: y = 16'h1ff;
			16'h118a: y = 16'h1ff;
			16'h118b: y = 16'h1ff;
			16'h118c: y = 16'h1ff;
			16'h118d: y = 16'h1ff;
			16'h118e: y = 16'h1ff;
			16'h118f: y = 16'h1ff;
			16'h1190: y = 16'h1ff;
			16'h1191: y = 16'h1ff;
			16'h1192: y = 16'h1ff;
			16'h1193: y = 16'h1ff;
			16'h1194: y = 16'h1ff;
			16'h1195: y = 16'h1ff;
			16'h1196: y = 16'h1ff;
			16'h1197: y = 16'h1ff;
			16'h1198: y = 16'h1ff;
			16'h1199: y = 16'h1ff;
			16'h119a: y = 16'h1ff;
			16'h119b: y = 16'h1ff;
			16'h119c: y = 16'h1ff;
			16'h119d: y = 16'h1ff;
			16'h119e: y = 16'h1ff;
			16'h119f: y = 16'h1ff;
			16'h11a0: y = 16'h1ff;
			16'h11a1: y = 16'h1ff;
			16'h11a2: y = 16'h1ff;
			16'h11a3: y = 16'h1ff;
			16'h11a4: y = 16'h1ff;
			16'h11a5: y = 16'h1ff;
			16'h11a6: y = 16'h1ff;
			16'h11a7: y = 16'h1ff;
			16'h11a8: y = 16'h1ff;
			16'h11a9: y = 16'h1ff;
			16'h11aa: y = 16'h1ff;
			16'h11ab: y = 16'h1ff;
			16'h11ac: y = 16'h1ff;
			16'h11ad: y = 16'h1ff;
			16'h11ae: y = 16'h1ff;
			16'h11af: y = 16'h1ff;
			16'h11b0: y = 16'h1ff;
			16'h11b1: y = 16'h1ff;
			16'h11b2: y = 16'h1ff;
			16'h11b3: y = 16'h1ff;
			16'h11b4: y = 16'h1ff;
			16'h11b5: y = 16'h1ff;
			16'h11b6: y = 16'h1ff;
			16'h11b7: y = 16'h1ff;
			16'h11b8: y = 16'h1ff;
			16'h11b9: y = 16'h1ff;
			16'h11ba: y = 16'h1ff;
			16'h11bb: y = 16'h1ff;
			16'h11bc: y = 16'h1ff;
			16'h11bd: y = 16'h1ff;
			16'h11be: y = 16'h1ff;
			16'h11bf: y = 16'h1ff;
			16'h11c0: y = 16'h1ff;
			16'h11c1: y = 16'h1ff;
			16'h11c2: y = 16'h1ff;
			16'h11c3: y = 16'h1ff;
			16'h11c4: y = 16'h1ff;
			16'h11c5: y = 16'h1ff;
			16'h11c6: y = 16'h1ff;
			16'h11c7: y = 16'h1ff;
			16'h11c8: y = 16'h1ff;
			16'h11c9: y = 16'h1ff;
			16'h11ca: y = 16'h1ff;
			16'h11cb: y = 16'h1ff;
			16'h11cc: y = 16'h1ff;
			16'h11cd: y = 16'h1ff;
			16'h11ce: y = 16'h1ff;
			16'h11cf: y = 16'h1ff;
			16'h11d0: y = 16'h1ff;
			16'h11d1: y = 16'h1ff;
			16'h11d2: y = 16'h1ff;
			16'h11d3: y = 16'h1ff;
			16'h11d4: y = 16'h1ff;
			16'h11d5: y = 16'h1ff;
			16'h11d6: y = 16'h1ff;
			16'h11d7: y = 16'h1ff;
			16'h11d8: y = 16'h1ff;
			16'h11d9: y = 16'h1ff;
			16'h11da: y = 16'h1ff;
			16'h11db: y = 16'h1ff;
			16'h11dc: y = 16'h1ff;
			16'h11dd: y = 16'h1ff;
			16'h11de: y = 16'h1ff;
			16'h11df: y = 16'h1ff;
			16'h11e0: y = 16'h1ff;
			16'h11e1: y = 16'h1ff;
			16'h11e2: y = 16'h1ff;
			16'h11e3: y = 16'h1ff;
			16'h11e4: y = 16'h1ff;
			16'h11e5: y = 16'h1ff;
			16'h11e6: y = 16'h1ff;
			16'h11e7: y = 16'h1ff;
			16'h11e8: y = 16'h1ff;
			16'h11e9: y = 16'h1ff;
			16'h11ea: y = 16'h1ff;
			16'h11eb: y = 16'h1ff;
			16'h11ec: y = 16'h1ff;
			16'h11ed: y = 16'h1ff;
			16'h11ee: y = 16'h1ff;
			16'h11ef: y = 16'h1ff;
			16'h11f0: y = 16'h1ff;
			16'h11f1: y = 16'h1ff;
			16'h11f2: y = 16'h1ff;
			16'h11f3: y = 16'h1ff;
			16'h11f4: y = 16'h1ff;
			16'h11f5: y = 16'h1ff;
			16'h11f6: y = 16'h1ff;
			16'h11f7: y = 16'h1ff;
			16'h11f8: y = 16'h1ff;
			16'h11f9: y = 16'h1ff;
			16'h11fa: y = 16'h1ff;
			16'h11fb: y = 16'h1ff;
			16'h11fc: y = 16'h1ff;
			16'h11fd: y = 16'h1ff;
			16'h11fe: y = 16'h1ff;
			16'h11ff: y = 16'h1ff;
			16'h1200: y = 16'h1ff;
			16'h1201: y = 16'h1ff;
			16'h1202: y = 16'h1ff;
			16'h1203: y = 16'h1ff;
			16'h1204: y = 16'h1ff;
			16'h1205: y = 16'h1ff;
			16'h1206: y = 16'h1ff;
			16'h1207: y = 16'h1ff;
			16'h1208: y = 16'h1ff;
			16'h1209: y = 16'h1ff;
			16'h120a: y = 16'h1ff;
			16'h120b: y = 16'h1ff;
			16'h120c: y = 16'h1ff;
			16'h120d: y = 16'h1ff;
			16'h120e: y = 16'h1ff;
			16'h120f: y = 16'h1ff;
			16'h1210: y = 16'h1ff;
			16'h1211: y = 16'h1ff;
			16'h1212: y = 16'h1ff;
			16'h1213: y = 16'h1ff;
			16'h1214: y = 16'h1ff;
			16'h1215: y = 16'h1ff;
			16'h1216: y = 16'h1ff;
			16'h1217: y = 16'h1ff;
			16'h1218: y = 16'h1ff;
			16'h1219: y = 16'h1ff;
			16'h121a: y = 16'h1ff;
			16'h121b: y = 16'h1ff;
			16'h121c: y = 16'h1ff;
			16'h121d: y = 16'h1ff;
			16'h121e: y = 16'h1ff;
			16'h121f: y = 16'h1ff;
			16'h1220: y = 16'h1ff;
			16'h1221: y = 16'h1ff;
			16'h1222: y = 16'h1ff;
			16'h1223: y = 16'h1ff;
			16'h1224: y = 16'h1ff;
			16'h1225: y = 16'h1ff;
			16'h1226: y = 16'h1ff;
			16'h1227: y = 16'h1ff;
			16'h1228: y = 16'h1ff;
			16'h1229: y = 16'h1ff;
			16'h122a: y = 16'h1ff;
			16'h122b: y = 16'h1ff;
			16'h122c: y = 16'h1ff;
			16'h122d: y = 16'h1ff;
			16'h122e: y = 16'h1ff;
			16'h122f: y = 16'h1ff;
			16'h1230: y = 16'h1ff;
			16'h1231: y = 16'h1ff;
			16'h1232: y = 16'h1ff;
			16'h1233: y = 16'h1ff;
			16'h1234: y = 16'h1ff;
			16'h1235: y = 16'h1ff;
			16'h1236: y = 16'h1ff;
			16'h1237: y = 16'h1ff;
			16'h1238: y = 16'h1ff;
			16'h1239: y = 16'h1ff;
			16'h123a: y = 16'h1ff;
			16'h123b: y = 16'h1ff;
			16'h123c: y = 16'h1ff;
			16'h123d: y = 16'h1ff;
			16'h123e: y = 16'h1ff;
			16'h123f: y = 16'h1ff;
			16'h1240: y = 16'h1ff;
			16'h1241: y = 16'h1ff;
			16'h1242: y = 16'h1ff;
			16'h1243: y = 16'h1ff;
			16'h1244: y = 16'h1ff;
			16'h1245: y = 16'h1ff;
			16'h1246: y = 16'h1ff;
			16'h1247: y = 16'h1ff;
			16'h1248: y = 16'h1ff;
			16'h1249: y = 16'h1ff;
			16'h124a: y = 16'h1ff;
			16'h124b: y = 16'h1ff;
			16'h124c: y = 16'h1ff;
			16'h124d: y = 16'h1ff;
			16'h124e: y = 16'h1ff;
			16'h124f: y = 16'h1ff;
			16'h1250: y = 16'h1ff;
			16'h1251: y = 16'h1ff;
			16'h1252: y = 16'h1ff;
			16'h1253: y = 16'h1ff;
			16'h1254: y = 16'h1ff;
			16'h1255: y = 16'h1ff;
			16'h1256: y = 16'h1ff;
			16'h1257: y = 16'h1ff;
			16'h1258: y = 16'h1ff;
			16'h1259: y = 16'h1ff;
			16'h125a: y = 16'h1ff;
			16'h125b: y = 16'h1ff;
			16'h125c: y = 16'h1ff;
			16'h125d: y = 16'h1ff;
			16'h125e: y = 16'h1ff;
			16'h125f: y = 16'h1ff;
			16'h1260: y = 16'h1ff;
			16'h1261: y = 16'h1ff;
			16'h1262: y = 16'h1ff;
			16'h1263: y = 16'h1ff;
			16'h1264: y = 16'h1ff;
			16'h1265: y = 16'h1ff;
			16'h1266: y = 16'h1ff;
			16'h1267: y = 16'h1ff;
			16'h1268: y = 16'h1ff;
			16'h1269: y = 16'h1ff;
			16'h126a: y = 16'h1ff;
			16'h126b: y = 16'h1ff;
			16'h126c: y = 16'h1ff;
			16'h126d: y = 16'h1ff;
			16'h126e: y = 16'h1ff;
			16'h126f: y = 16'h1ff;
			16'h1270: y = 16'h1ff;
			16'h1271: y = 16'h1ff;
			16'h1272: y = 16'h1ff;
			16'h1273: y = 16'h1ff;
			16'h1274: y = 16'h1ff;
			16'h1275: y = 16'h1ff;
			16'h1276: y = 16'h1ff;
			16'h1277: y = 16'h1ff;
			16'h1278: y = 16'h1ff;
			16'h1279: y = 16'h1ff;
			16'h127a: y = 16'h1ff;
			16'h127b: y = 16'h1ff;
			16'h127c: y = 16'h1ff;
			16'h127d: y = 16'h1ff;
			16'h127e: y = 16'h1ff;
			16'h127f: y = 16'h1ff;
			16'h1280: y = 16'h1ff;
			16'h1281: y = 16'h1ff;
			16'h1282: y = 16'h1ff;
			16'h1283: y = 16'h1ff;
			16'h1284: y = 16'h1ff;
			16'h1285: y = 16'h1ff;
			16'h1286: y = 16'h1ff;
			16'h1287: y = 16'h1ff;
			16'h1288: y = 16'h1ff;
			16'h1289: y = 16'h1ff;
			16'h128a: y = 16'h1ff;
			16'h128b: y = 16'h1ff;
			16'h128c: y = 16'h1ff;
			16'h128d: y = 16'h1ff;
			16'h128e: y = 16'h1ff;
			16'h128f: y = 16'h1ff;
			16'h1290: y = 16'h1ff;
			16'h1291: y = 16'h1ff;
			16'h1292: y = 16'h1ff;
			16'h1293: y = 16'h1ff;
			16'h1294: y = 16'h1ff;
			16'h1295: y = 16'h1ff;
			16'h1296: y = 16'h1ff;
			16'h1297: y = 16'h1ff;
			16'h1298: y = 16'h1ff;
			16'h1299: y = 16'h1ff;
			16'h129a: y = 16'h1ff;
			16'h129b: y = 16'h1ff;
			16'h129c: y = 16'h1ff;
			16'h129d: y = 16'h1ff;
			16'h129e: y = 16'h1ff;
			16'h129f: y = 16'h1ff;
			16'h12a0: y = 16'h1ff;
			16'h12a1: y = 16'h1ff;
			16'h12a2: y = 16'h1ff;
			16'h12a3: y = 16'h1ff;
			16'h12a4: y = 16'h1ff;
			16'h12a5: y = 16'h1ff;
			16'h12a6: y = 16'h1ff;
			16'h12a7: y = 16'h1ff;
			16'h12a8: y = 16'h1ff;
			16'h12a9: y = 16'h1ff;
			16'h12aa: y = 16'h1ff;
			16'h12ab: y = 16'h1ff;
			16'h12ac: y = 16'h1ff;
			16'h12ad: y = 16'h1ff;
			16'h12ae: y = 16'h1ff;
			16'h12af: y = 16'h1ff;
			16'h12b0: y = 16'h1ff;
			16'h12b1: y = 16'h1ff;
			16'h12b2: y = 16'h1ff;
			16'h12b3: y = 16'h1ff;
			16'h12b4: y = 16'h1ff;
			16'h12b5: y = 16'h1ff;
			16'h12b6: y = 16'h1ff;
			16'h12b7: y = 16'h1ff;
			16'h12b8: y = 16'h1ff;
			16'h12b9: y = 16'h1ff;
			16'h12ba: y = 16'h1ff;
			16'h12bb: y = 16'h1ff;
			16'h12bc: y = 16'h1ff;
			16'h12bd: y = 16'h1ff;
			16'h12be: y = 16'h1ff;
			16'h12bf: y = 16'h1ff;
			16'h12c0: y = 16'h1ff;
			16'h12c1: y = 16'h1ff;
			16'h12c2: y = 16'h1ff;
			16'h12c3: y = 16'h1ff;
			16'h12c4: y = 16'h1ff;
			16'h12c5: y = 16'h1ff;
			16'h12c6: y = 16'h1ff;
			16'h12c7: y = 16'h1ff;
			16'h12c8: y = 16'h1ff;
			16'h12c9: y = 16'h1ff;
			16'h12ca: y = 16'h1ff;
			16'h12cb: y = 16'h1ff;
			16'h12cc: y = 16'h1ff;
			16'h12cd: y = 16'h1ff;
			16'h12ce: y = 16'h1ff;
			16'h12cf: y = 16'h1ff;
			16'h12d0: y = 16'h1ff;
			16'h12d1: y = 16'h1ff;
			16'h12d2: y = 16'h1ff;
			16'h12d3: y = 16'h1ff;
			16'h12d4: y = 16'h1ff;
			16'h12d5: y = 16'h1ff;
			16'h12d6: y = 16'h1ff;
			16'h12d7: y = 16'h1ff;
			16'h12d8: y = 16'h1ff;
			16'h12d9: y = 16'h1ff;
			16'h12da: y = 16'h1ff;
			16'h12db: y = 16'h1ff;
			16'h12dc: y = 16'h1ff;
			16'h12dd: y = 16'h1ff;
			16'h12de: y = 16'h1ff;
			16'h12df: y = 16'h1ff;
			16'h12e0: y = 16'h1ff;
			16'h12e1: y = 16'h1ff;
			16'h12e2: y = 16'h1ff;
			16'h12e3: y = 16'h1ff;
			16'h12e4: y = 16'h1ff;
			16'h12e5: y = 16'h1ff;
			16'h12e6: y = 16'h1ff;
			16'h12e7: y = 16'h1ff;
			16'h12e8: y = 16'h1ff;
			16'h12e9: y = 16'h1ff;
			16'h12ea: y = 16'h1ff;
			16'h12eb: y = 16'h1ff;
			16'h12ec: y = 16'h1ff;
			16'h12ed: y = 16'h1ff;
			16'h12ee: y = 16'h1ff;
			16'h12ef: y = 16'h1ff;
			16'h12f0: y = 16'h1ff;
			16'h12f1: y = 16'h1ff;
			16'h12f2: y = 16'h1ff;
			16'h12f3: y = 16'h1ff;
			16'h12f4: y = 16'h1ff;
			16'h12f5: y = 16'h1ff;
			16'h12f6: y = 16'h1ff;
			16'h12f7: y = 16'h1ff;
			16'h12f8: y = 16'h1ff;
			16'h12f9: y = 16'h1ff;
			16'h12fa: y = 16'h1ff;
			16'h12fb: y = 16'h1ff;
			16'h12fc: y = 16'h1ff;
			16'h12fd: y = 16'h1ff;
			16'h12fe: y = 16'h1ff;
			16'h12ff: y = 16'h1ff;
			16'h1300: y = 16'h1ff;
			16'h1301: y = 16'h1ff;
			16'h1302: y = 16'h1ff;
			16'h1303: y = 16'h1ff;
			16'h1304: y = 16'h1ff;
			16'h1305: y = 16'h1ff;
			16'h1306: y = 16'h1ff;
			16'h1307: y = 16'h1ff;
			16'h1308: y = 16'h1ff;
			16'h1309: y = 16'h1ff;
			16'h130a: y = 16'h1ff;
			16'h130b: y = 16'h1ff;
			16'h130c: y = 16'h1ff;
			16'h130d: y = 16'h1ff;
			16'h130e: y = 16'h1ff;
			16'h130f: y = 16'h1ff;
			16'h1310: y = 16'h1ff;
			16'h1311: y = 16'h1ff;
			16'h1312: y = 16'h1ff;
			16'h1313: y = 16'h1ff;
			16'h1314: y = 16'h1ff;
			16'h1315: y = 16'h1ff;
			16'h1316: y = 16'h1ff;
			16'h1317: y = 16'h1ff;
			16'h1318: y = 16'h1ff;
			16'h1319: y = 16'h1ff;
			16'h131a: y = 16'h1ff;
			16'h131b: y = 16'h1ff;
			16'h131c: y = 16'h1ff;
			16'h131d: y = 16'h1ff;
			16'h131e: y = 16'h1ff;
			16'h131f: y = 16'h1ff;
			16'h1320: y = 16'h1ff;
			16'h1321: y = 16'h1ff;
			16'h1322: y = 16'h1ff;
			16'h1323: y = 16'h1ff;
			16'h1324: y = 16'h1ff;
			16'h1325: y = 16'h1ff;
			16'h1326: y = 16'h1ff;
			16'h1327: y = 16'h1ff;
			16'h1328: y = 16'h1ff;
			16'h1329: y = 16'h1ff;
			16'h132a: y = 16'h1ff;
			16'h132b: y = 16'h1ff;
			16'h132c: y = 16'h1ff;
			16'h132d: y = 16'h1ff;
			16'h132e: y = 16'h1ff;
			16'h132f: y = 16'h1ff;
			16'h1330: y = 16'h1ff;
			16'h1331: y = 16'h1ff;
			16'h1332: y = 16'h1ff;
			16'h1333: y = 16'h1ff;
			16'h1334: y = 16'h1ff;
			16'h1335: y = 16'h1ff;
			16'h1336: y = 16'h1ff;
			16'h1337: y = 16'h1ff;
			16'h1338: y = 16'h1ff;
			16'h1339: y = 16'h1ff;
			16'h133a: y = 16'h1ff;
			16'h133b: y = 16'h1ff;
			16'h133c: y = 16'h1ff;
			16'h133d: y = 16'h1ff;
			16'h133e: y = 16'h1ff;
			16'h133f: y = 16'h1ff;
			16'h1340: y = 16'h1ff;
			16'h1341: y = 16'h1ff;
			16'h1342: y = 16'h1ff;
			16'h1343: y = 16'h1ff;
			16'h1344: y = 16'h1ff;
			16'h1345: y = 16'h1ff;
			16'h1346: y = 16'h1ff;
			16'h1347: y = 16'h1ff;
			16'h1348: y = 16'h1ff;
			16'h1349: y = 16'h1ff;
			16'h134a: y = 16'h1ff;
			16'h134b: y = 16'h1ff;
			16'h134c: y = 16'h1ff;
			16'h134d: y = 16'h1ff;
			16'h134e: y = 16'h1ff;
			16'h134f: y = 16'h1ff;
			16'h1350: y = 16'h1ff;
			16'h1351: y = 16'h1ff;
			16'h1352: y = 16'h1ff;
			16'h1353: y = 16'h1ff;
			16'h1354: y = 16'h1ff;
			16'h1355: y = 16'h1ff;
			16'h1356: y = 16'h1ff;
			16'h1357: y = 16'h1ff;
			16'h1358: y = 16'h1ff;
			16'h1359: y = 16'h1ff;
			16'h135a: y = 16'h1ff;
			16'h135b: y = 16'h1ff;
			16'h135c: y = 16'h1ff;
			16'h135d: y = 16'h1ff;
			16'h135e: y = 16'h1ff;
			16'h135f: y = 16'h1ff;
			16'h1360: y = 16'h1ff;
			16'h1361: y = 16'h1ff;
			16'h1362: y = 16'h1ff;
			16'h1363: y = 16'h1ff;
			16'h1364: y = 16'h1ff;
			16'h1365: y = 16'h1ff;
			16'h1366: y = 16'h1ff;
			16'h1367: y = 16'h1ff;
			16'h1368: y = 16'h1ff;
			16'h1369: y = 16'h1ff;
			16'h136a: y = 16'h1ff;
			16'h136b: y = 16'h1ff;
			16'h136c: y = 16'h1ff;
			16'h136d: y = 16'h1ff;
			16'h136e: y = 16'h1ff;
			16'h136f: y = 16'h1ff;
			16'h1370: y = 16'h1ff;
			16'h1371: y = 16'h1ff;
			16'h1372: y = 16'h1ff;
			16'h1373: y = 16'h1ff;
			16'h1374: y = 16'h1ff;
			16'h1375: y = 16'h1ff;
			16'h1376: y = 16'h1ff;
			16'h1377: y = 16'h1ff;
			16'h1378: y = 16'h1ff;
			16'h1379: y = 16'h1ff;
			16'h137a: y = 16'h1ff;
			16'h137b: y = 16'h1ff;
			16'h137c: y = 16'h1ff;
			16'h137d: y = 16'h1ff;
			16'h137e: y = 16'h1ff;
			16'h137f: y = 16'h1ff;
			16'h1380: y = 16'h1ff;
			16'h1381: y = 16'h1ff;
			16'h1382: y = 16'h1ff;
			16'h1383: y = 16'h1ff;
			16'h1384: y = 16'h1ff;
			16'h1385: y = 16'h1ff;
			16'h1386: y = 16'h1ff;
			16'h1387: y = 16'h1ff;
			16'h1388: y = 16'h1ff;
			16'h1389: y = 16'h1ff;
			16'h138a: y = 16'h1ff;
			16'h138b: y = 16'h1ff;
			16'h138c: y = 16'h1ff;
			16'h138d: y = 16'h1ff;
			16'h138e: y = 16'h1ff;
			16'h138f: y = 16'h1ff;
			16'h1390: y = 16'h1ff;
			16'h1391: y = 16'h1ff;
			16'h1392: y = 16'h1ff;
			16'h1393: y = 16'h1ff;
			16'h1394: y = 16'h1ff;
			16'h1395: y = 16'h1ff;
			16'h1396: y = 16'h1ff;
			16'h1397: y = 16'h1ff;
			16'h1398: y = 16'h1ff;
			16'h1399: y = 16'h1ff;
			16'h139a: y = 16'h1ff;
			16'h139b: y = 16'h1ff;
			16'h139c: y = 16'h1ff;
			16'h139d: y = 16'h1ff;
			16'h139e: y = 16'h1ff;
			16'h139f: y = 16'h1ff;
			16'h13a0: y = 16'h1ff;
			16'h13a1: y = 16'h1ff;
			16'h13a2: y = 16'h1ff;
			16'h13a3: y = 16'h1ff;
			16'h13a4: y = 16'h1ff;
			16'h13a5: y = 16'h1ff;
			16'h13a6: y = 16'h1ff;
			16'h13a7: y = 16'h1ff;
			16'h13a8: y = 16'h1ff;
			16'h13a9: y = 16'h1ff;
			16'h13aa: y = 16'h1ff;
			16'h13ab: y = 16'h1ff;
			16'h13ac: y = 16'h1ff;
			16'h13ad: y = 16'h1ff;
			16'h13ae: y = 16'h1ff;
			16'h13af: y = 16'h1ff;
			16'h13b0: y = 16'h1ff;
			16'h13b1: y = 16'h1ff;
			16'h13b2: y = 16'h1ff;
			16'h13b3: y = 16'h1ff;
			16'h13b4: y = 16'h1ff;
			16'h13b5: y = 16'h1ff;
			16'h13b6: y = 16'h1ff;
			16'h13b7: y = 16'h1ff;
			16'h13b8: y = 16'h1ff;
			16'h13b9: y = 16'h1ff;
			16'h13ba: y = 16'h1ff;
			16'h13bb: y = 16'h1ff;
			16'h13bc: y = 16'h1ff;
			16'h13bd: y = 16'h1ff;
			16'h13be: y = 16'h1ff;
			16'h13bf: y = 16'h1ff;
			16'h13c0: y = 16'h1ff;
			16'h13c1: y = 16'h1ff;
			16'h13c2: y = 16'h1ff;
			16'h13c3: y = 16'h1ff;
			16'h13c4: y = 16'h1ff;
			16'h13c5: y = 16'h1ff;
			16'h13c6: y = 16'h1ff;
			16'h13c7: y = 16'h1ff;
			16'h13c8: y = 16'h1ff;
			16'h13c9: y = 16'h1ff;
			16'h13ca: y = 16'h1ff;
			16'h13cb: y = 16'h1ff;
			16'h13cc: y = 16'h1ff;
			16'h13cd: y = 16'h1ff;
			16'h13ce: y = 16'h1ff;
			16'h13cf: y = 16'h1ff;
			16'h13d0: y = 16'h1ff;
			16'h13d1: y = 16'h1ff;
			16'h13d2: y = 16'h1ff;
			16'h13d3: y = 16'h1ff;
			16'h13d4: y = 16'h1ff;
			16'h13d5: y = 16'h1ff;
			16'h13d6: y = 16'h1ff;
			16'h13d7: y = 16'h1ff;
			16'h13d8: y = 16'h1ff;
			16'h13d9: y = 16'h1ff;
			16'h13da: y = 16'h1ff;
			16'h13db: y = 16'h1ff;
			16'h13dc: y = 16'h1ff;
			16'h13dd: y = 16'h1ff;
			16'h13de: y = 16'h1ff;
			16'h13df: y = 16'h1ff;
			16'h13e0: y = 16'h1ff;
			16'h13e1: y = 16'h1ff;
			16'h13e2: y = 16'h1ff;
			16'h13e3: y = 16'h1ff;
			16'h13e4: y = 16'h1ff;
			16'h13e5: y = 16'h1ff;
			16'h13e6: y = 16'h1ff;
			16'h13e7: y = 16'h1ff;
			16'h13e8: y = 16'h1ff;
			16'h13e9: y = 16'h1ff;
			16'h13ea: y = 16'h1ff;
			16'h13eb: y = 16'h1ff;
			16'h13ec: y = 16'h1ff;
			16'h13ed: y = 16'h1ff;
			16'h13ee: y = 16'h1ff;
			16'h13ef: y = 16'h1ff;
			16'h13f0: y = 16'h1ff;
			16'h13f1: y = 16'h1ff;
			16'h13f2: y = 16'h1ff;
			16'h13f3: y = 16'h1ff;
			16'h13f4: y = 16'h1ff;
			16'h13f5: y = 16'h1ff;
			16'h13f6: y = 16'h1ff;
			16'h13f7: y = 16'h1ff;
			16'h13f8: y = 16'h1ff;
			16'h13f9: y = 16'h1ff;
			16'h13fa: y = 16'h1ff;
			16'h13fb: y = 16'h1ff;
			16'h13fc: y = 16'h1ff;
			16'h13fd: y = 16'h1ff;
			16'h13fe: y = 16'h1ff;
			16'h13ff: y = 16'h1ff;
			16'h1400: y = 16'h1ff;
			16'h1401: y = 16'h1ff;
			16'h1402: y = 16'h1ff;
			16'h1403: y = 16'h1ff;
			16'h1404: y = 16'h1ff;
			16'h1405: y = 16'h1ff;
			16'h1406: y = 16'h1ff;
			16'h1407: y = 16'h1ff;
			16'h1408: y = 16'h1ff;
			16'h1409: y = 16'h1ff;
			16'h140a: y = 16'h1ff;
			16'h140b: y = 16'h1ff;
			16'h140c: y = 16'h1ff;
			16'h140d: y = 16'h1ff;
			16'h140e: y = 16'h1ff;
			16'h140f: y = 16'h1ff;
			16'h1410: y = 16'h1ff;
			16'h1411: y = 16'h1ff;
			16'h1412: y = 16'h1ff;
			16'h1413: y = 16'h1ff;
			16'h1414: y = 16'h1ff;
			16'h1415: y = 16'h1ff;
			16'h1416: y = 16'h1ff;
			16'h1417: y = 16'h1ff;
			16'h1418: y = 16'h1ff;
			16'h1419: y = 16'h1ff;
			16'h141a: y = 16'h1ff;
			16'h141b: y = 16'h1ff;
			16'h141c: y = 16'h1ff;
			16'h141d: y = 16'h1ff;
			16'h141e: y = 16'h1ff;
			16'h141f: y = 16'h1ff;
			16'h1420: y = 16'h1ff;
			16'h1421: y = 16'h1ff;
			16'h1422: y = 16'h1ff;
			16'h1423: y = 16'h1ff;
			16'h1424: y = 16'h1ff;
			16'h1425: y = 16'h1ff;
			16'h1426: y = 16'h1ff;
			16'h1427: y = 16'h1ff;
			16'h1428: y = 16'h1ff;
			16'h1429: y = 16'h1ff;
			16'h142a: y = 16'h1ff;
			16'h142b: y = 16'h1ff;
			16'h142c: y = 16'h1ff;
			16'h142d: y = 16'h1ff;
			16'h142e: y = 16'h1ff;
			16'h142f: y = 16'h1ff;
			16'h1430: y = 16'h1ff;
			16'h1431: y = 16'h1ff;
			16'h1432: y = 16'h1ff;
			16'h1433: y = 16'h1ff;
			16'h1434: y = 16'h1ff;
			16'h1435: y = 16'h1ff;
			16'h1436: y = 16'h1ff;
			16'h1437: y = 16'h1ff;
			16'h1438: y = 16'h1ff;
			16'h1439: y = 16'h1ff;
			16'h143a: y = 16'h1ff;
			16'h143b: y = 16'h1ff;
			16'h143c: y = 16'h1ff;
			16'h143d: y = 16'h1ff;
			16'h143e: y = 16'h1ff;
			16'h143f: y = 16'h1ff;
			16'h1440: y = 16'h1ff;
			16'h1441: y = 16'h1ff;
			16'h1442: y = 16'h1ff;
			16'h1443: y = 16'h1ff;
			16'h1444: y = 16'h1ff;
			16'h1445: y = 16'h1ff;
			16'h1446: y = 16'h1ff;
			16'h1447: y = 16'h1ff;
			16'h1448: y = 16'h1ff;
			16'h1449: y = 16'h1ff;
			16'h144a: y = 16'h1ff;
			16'h144b: y = 16'h1ff;
			16'h144c: y = 16'h1ff;
			16'h144d: y = 16'h1ff;
			16'h144e: y = 16'h1ff;
			16'h144f: y = 16'h1ff;
			16'h1450: y = 16'h1ff;
			16'h1451: y = 16'h1ff;
			16'h1452: y = 16'h1ff;
			16'h1453: y = 16'h1ff;
			16'h1454: y = 16'h1ff;
			16'h1455: y = 16'h1ff;
			16'h1456: y = 16'h1ff;
			16'h1457: y = 16'h1ff;
			16'h1458: y = 16'h1ff;
			16'h1459: y = 16'h1ff;
			16'h145a: y = 16'h1ff;
			16'h145b: y = 16'h1ff;
			16'h145c: y = 16'h1ff;
			16'h145d: y = 16'h1ff;
			16'h145e: y = 16'h1ff;
			16'h145f: y = 16'h1ff;
			16'h1460: y = 16'h1ff;
			16'h1461: y = 16'h1ff;
			16'h1462: y = 16'h1ff;
			16'h1463: y = 16'h1ff;
			16'h1464: y = 16'h1ff;
			16'h1465: y = 16'h1ff;
			16'h1466: y = 16'h1ff;
			16'h1467: y = 16'h1ff;
			16'h1468: y = 16'h1ff;
			16'h1469: y = 16'h1ff;
			16'h146a: y = 16'h1ff;
			16'h146b: y = 16'h1ff;
			16'h146c: y = 16'h1ff;
			16'h146d: y = 16'h1ff;
			16'h146e: y = 16'h1ff;
			16'h146f: y = 16'h1ff;
			16'h1470: y = 16'h1ff;
			16'h1471: y = 16'h1ff;
			16'h1472: y = 16'h1ff;
			16'h1473: y = 16'h1ff;
			16'h1474: y = 16'h1ff;
			16'h1475: y = 16'h1ff;
			16'h1476: y = 16'h1ff;
			16'h1477: y = 16'h1ff;
			16'h1478: y = 16'h1ff;
			16'h1479: y = 16'h1ff;
			16'h147a: y = 16'h1ff;
			16'h147b: y = 16'h1ff;
			16'h147c: y = 16'h1ff;
			16'h147d: y = 16'h1ff;
			16'h147e: y = 16'h1ff;
			16'h147f: y = 16'h1ff;
			16'h1480: y = 16'h1ff;
			16'h1481: y = 16'h1ff;
			16'h1482: y = 16'h1ff;
			16'h1483: y = 16'h1ff;
			16'h1484: y = 16'h1ff;
			16'h1485: y = 16'h1ff;
			16'h1486: y = 16'h1ff;
			16'h1487: y = 16'h1ff;
			16'h1488: y = 16'h1ff;
			16'h1489: y = 16'h1ff;
			16'h148a: y = 16'h1ff;
			16'h148b: y = 16'h1ff;
			16'h148c: y = 16'h1ff;
			16'h148d: y = 16'h1ff;
			16'h148e: y = 16'h1ff;
			16'h148f: y = 16'h1ff;
			16'h1490: y = 16'h1ff;
			16'h1491: y = 16'h1ff;
			16'h1492: y = 16'h1ff;
			16'h1493: y = 16'h1ff;
			16'h1494: y = 16'h1ff;
			16'h1495: y = 16'h1ff;
			16'h1496: y = 16'h1ff;
			16'h1497: y = 16'h1ff;
			16'h1498: y = 16'h1ff;
			16'h1499: y = 16'h1ff;
			16'h149a: y = 16'h1ff;
			16'h149b: y = 16'h1ff;
			16'h149c: y = 16'h1ff;
			16'h149d: y = 16'h1ff;
			16'h149e: y = 16'h1ff;
			16'h149f: y = 16'h1ff;
			16'h14a0: y = 16'h1ff;
			16'h14a1: y = 16'h1ff;
			16'h14a2: y = 16'h1ff;
			16'h14a3: y = 16'h1ff;
			16'h14a4: y = 16'h1ff;
			16'h14a5: y = 16'h1ff;
			16'h14a6: y = 16'h1ff;
			16'h14a7: y = 16'h1ff;
			16'h14a8: y = 16'h1ff;
			16'h14a9: y = 16'h1ff;
			16'h14aa: y = 16'h1ff;
			16'h14ab: y = 16'h1ff;
			16'h14ac: y = 16'h1ff;
			16'h14ad: y = 16'h1ff;
			16'h14ae: y = 16'h1ff;
			16'h14af: y = 16'h1ff;
			16'h14b0: y = 16'h1ff;
			16'h14b1: y = 16'h1ff;
			16'h14b2: y = 16'h1ff;
			16'h14b3: y = 16'h1ff;
			16'h14b4: y = 16'h1ff;
			16'h14b5: y = 16'h1ff;
			16'h14b6: y = 16'h1ff;
			16'h14b7: y = 16'h1ff;
			16'h14b8: y = 16'h1ff;
			16'h14b9: y = 16'h1ff;
			16'h14ba: y = 16'h1ff;
			16'h14bb: y = 16'h1ff;
			16'h14bc: y = 16'h1ff;
			16'h14bd: y = 16'h1ff;
			16'h14be: y = 16'h1ff;
			16'h14bf: y = 16'h1ff;
			16'h14c0: y = 16'h1ff;
			16'h14c1: y = 16'h1ff;
			16'h14c2: y = 16'h1ff;
			16'h14c3: y = 16'h1ff;
			16'h14c4: y = 16'h1ff;
			16'h14c5: y = 16'h1ff;
			16'h14c6: y = 16'h1ff;
			16'h14c7: y = 16'h1ff;
			16'h14c8: y = 16'h1ff;
			16'h14c9: y = 16'h1ff;
			16'h14ca: y = 16'h1ff;
			16'h14cb: y = 16'h1ff;
			16'h14cc: y = 16'h1ff;
			16'h14cd: y = 16'h1ff;
			16'h14ce: y = 16'h1ff;
			16'h14cf: y = 16'h1ff;
			16'h14d0: y = 16'h1ff;
			16'h14d1: y = 16'h1ff;
			16'h14d2: y = 16'h1ff;
			16'h14d3: y = 16'h1ff;
			16'h14d4: y = 16'h1ff;
			16'h14d5: y = 16'h1ff;
			16'h14d6: y = 16'h1ff;
			16'h14d7: y = 16'h1ff;
			16'h14d8: y = 16'h1ff;
			16'h14d9: y = 16'h1ff;
			16'h14da: y = 16'h1ff;
			16'h14db: y = 16'h1ff;
			16'h14dc: y = 16'h1ff;
			16'h14dd: y = 16'h1ff;
			16'h14de: y = 16'h1ff;
			16'h14df: y = 16'h1ff;
			16'h14e0: y = 16'h1ff;
			16'h14e1: y = 16'h1ff;
			16'h14e2: y = 16'h1ff;
			16'h14e3: y = 16'h1ff;
			16'h14e4: y = 16'h1ff;
			16'h14e5: y = 16'h1ff;
			16'h14e6: y = 16'h1ff;
			16'h14e7: y = 16'h1ff;
			16'h14e8: y = 16'h1ff;
			16'h14e9: y = 16'h1ff;
			16'h14ea: y = 16'h1ff;
			16'h14eb: y = 16'h1ff;
			16'h14ec: y = 16'h1ff;
			16'h14ed: y = 16'h1ff;
			16'h14ee: y = 16'h1ff;
			16'h14ef: y = 16'h1ff;
			16'h14f0: y = 16'h1ff;
			16'h14f1: y = 16'h1ff;
			16'h14f2: y = 16'h1ff;
			16'h14f3: y = 16'h1ff;
			16'h14f4: y = 16'h1ff;
			16'h14f5: y = 16'h1ff;
			16'h14f6: y = 16'h1ff;
			16'h14f7: y = 16'h1ff;
			16'h14f8: y = 16'h1ff;
			16'h14f9: y = 16'h1ff;
			16'h14fa: y = 16'h1ff;
			16'h14fb: y = 16'h1ff;
			16'h14fc: y = 16'h1ff;
			16'h14fd: y = 16'h1ff;
			16'h14fe: y = 16'h1ff;
			16'h14ff: y = 16'h1ff;
			16'h1500: y = 16'h1ff;
			16'h1501: y = 16'h1ff;
			16'h1502: y = 16'h1ff;
			16'h1503: y = 16'h1ff;
			16'h1504: y = 16'h1ff;
			16'h1505: y = 16'h1ff;
			16'h1506: y = 16'h1ff;
			16'h1507: y = 16'h1ff;
			16'h1508: y = 16'h1ff;
			16'h1509: y = 16'h1ff;
			16'h150a: y = 16'h1ff;
			16'h150b: y = 16'h1ff;
			16'h150c: y = 16'h1ff;
			16'h150d: y = 16'h1ff;
			16'h150e: y = 16'h1ff;
			16'h150f: y = 16'h1ff;
			16'h1510: y = 16'h1ff;
			16'h1511: y = 16'h1ff;
			16'h1512: y = 16'h1ff;
			16'h1513: y = 16'h1ff;
			16'h1514: y = 16'h1ff;
			16'h1515: y = 16'h1ff;
			16'h1516: y = 16'h1ff;
			16'h1517: y = 16'h1ff;
			16'h1518: y = 16'h1ff;
			16'h1519: y = 16'h1ff;
			16'h151a: y = 16'h1ff;
			16'h151b: y = 16'h1ff;
			16'h151c: y = 16'h1ff;
			16'h151d: y = 16'h1ff;
			16'h151e: y = 16'h1ff;
			16'h151f: y = 16'h1ff;
			16'h1520: y = 16'h1ff;
			16'h1521: y = 16'h1ff;
			16'h1522: y = 16'h1ff;
			16'h1523: y = 16'h1ff;
			16'h1524: y = 16'h1ff;
			16'h1525: y = 16'h1ff;
			16'h1526: y = 16'h1ff;
			16'h1527: y = 16'h1ff;
			16'h1528: y = 16'h1ff;
			16'h1529: y = 16'h1ff;
			16'h152a: y = 16'h1ff;
			16'h152b: y = 16'h1ff;
			16'h152c: y = 16'h1ff;
			16'h152d: y = 16'h1ff;
			16'h152e: y = 16'h1ff;
			16'h152f: y = 16'h1ff;
			16'h1530: y = 16'h1ff;
			16'h1531: y = 16'h1ff;
			16'h1532: y = 16'h1ff;
			16'h1533: y = 16'h1ff;
			16'h1534: y = 16'h1ff;
			16'h1535: y = 16'h1ff;
			16'h1536: y = 16'h1ff;
			16'h1537: y = 16'h1ff;
			16'h1538: y = 16'h1ff;
			16'h1539: y = 16'h1ff;
			16'h153a: y = 16'h1ff;
			16'h153b: y = 16'h1ff;
			16'h153c: y = 16'h1ff;
			16'h153d: y = 16'h1ff;
			16'h153e: y = 16'h1ff;
			16'h153f: y = 16'h1ff;
			16'h1540: y = 16'h1ff;
			16'h1541: y = 16'h1ff;
			16'h1542: y = 16'h1ff;
			16'h1543: y = 16'h1ff;
			16'h1544: y = 16'h1ff;
			16'h1545: y = 16'h1ff;
			16'h1546: y = 16'h1ff;
			16'h1547: y = 16'h1ff;
			16'h1548: y = 16'h1ff;
			16'h1549: y = 16'h1ff;
			16'h154a: y = 16'h1ff;
			16'h154b: y = 16'h1ff;
			16'h154c: y = 16'h1ff;
			16'h154d: y = 16'h1ff;
			16'h154e: y = 16'h1ff;
			16'h154f: y = 16'h1ff;
			16'h1550: y = 16'h1ff;
			16'h1551: y = 16'h1ff;
			16'h1552: y = 16'h1ff;
			16'h1553: y = 16'h1ff;
			16'h1554: y = 16'h1ff;
			16'h1555: y = 16'h1ff;
			16'h1556: y = 16'h1ff;
			16'h1557: y = 16'h1ff;
			16'h1558: y = 16'h1ff;
			16'h1559: y = 16'h1ff;
			16'h155a: y = 16'h1ff;
			16'h155b: y = 16'h1ff;
			16'h155c: y = 16'h1ff;
			16'h155d: y = 16'h1ff;
			16'h155e: y = 16'h1ff;
			16'h155f: y = 16'h1ff;
			16'h1560: y = 16'h1ff;
			16'h1561: y = 16'h1ff;
			16'h1562: y = 16'h1ff;
			16'h1563: y = 16'h1ff;
			16'h1564: y = 16'h1ff;
			16'h1565: y = 16'h1ff;
			16'h1566: y = 16'h1ff;
			16'h1567: y = 16'h1ff;
			16'h1568: y = 16'h1ff;
			16'h1569: y = 16'h1ff;
			16'h156a: y = 16'h1ff;
			16'h156b: y = 16'h1ff;
			16'h156c: y = 16'h1ff;
			16'h156d: y = 16'h1ff;
			16'h156e: y = 16'h1ff;
			16'h156f: y = 16'h1ff;
			16'h1570: y = 16'h1ff;
			16'h1571: y = 16'h1ff;
			16'h1572: y = 16'h1ff;
			16'h1573: y = 16'h1ff;
			16'h1574: y = 16'h1ff;
			16'h1575: y = 16'h1ff;
			16'h1576: y = 16'h1ff;
			16'h1577: y = 16'h1ff;
			16'h1578: y = 16'h1ff;
			16'h1579: y = 16'h1ff;
			16'h157a: y = 16'h1ff;
			16'h157b: y = 16'h1ff;
			16'h157c: y = 16'h1ff;
			16'h157d: y = 16'h1ff;
			16'h157e: y = 16'h1ff;
			16'h157f: y = 16'h1ff;
			16'h1580: y = 16'h1ff;
			16'h1581: y = 16'h1ff;
			16'h1582: y = 16'h1ff;
			16'h1583: y = 16'h1ff;
			16'h1584: y = 16'h1ff;
			16'h1585: y = 16'h1ff;
			16'h1586: y = 16'h1ff;
			16'h1587: y = 16'h1ff;
			16'h1588: y = 16'h1ff;
			16'h1589: y = 16'h1ff;
			16'h158a: y = 16'h1ff;
			16'h158b: y = 16'h1ff;
			16'h158c: y = 16'h1ff;
			16'h158d: y = 16'h1ff;
			16'h158e: y = 16'h1ff;
			16'h158f: y = 16'h1ff;
			16'h1590: y = 16'h1ff;
			16'h1591: y = 16'h1ff;
			16'h1592: y = 16'h1ff;
			16'h1593: y = 16'h1ff;
			16'h1594: y = 16'h1ff;
			16'h1595: y = 16'h1ff;
			16'h1596: y = 16'h1ff;
			16'h1597: y = 16'h1ff;
			16'h1598: y = 16'h1ff;
			16'h1599: y = 16'h1ff;
			16'h159a: y = 16'h1ff;
			16'h159b: y = 16'h1ff;
			16'h159c: y = 16'h1ff;
			16'h159d: y = 16'h1ff;
			16'h159e: y = 16'h1ff;
			16'h159f: y = 16'h1ff;
			16'h15a0: y = 16'h1ff;
			16'h15a1: y = 16'h1ff;
			16'h15a2: y = 16'h1ff;
			16'h15a3: y = 16'h1ff;
			16'h15a4: y = 16'h1ff;
			16'h15a5: y = 16'h1ff;
			16'h15a6: y = 16'h1ff;
			16'h15a7: y = 16'h1ff;
			16'h15a8: y = 16'h1ff;
			16'h15a9: y = 16'h1ff;
			16'h15aa: y = 16'h1ff;
			16'h15ab: y = 16'h1ff;
			16'h15ac: y = 16'h1ff;
			16'h15ad: y = 16'h1ff;
			16'h15ae: y = 16'h1ff;
			16'h15af: y = 16'h1ff;
			16'h15b0: y = 16'h1ff;
			16'h15b1: y = 16'h1ff;
			16'h15b2: y = 16'h1ff;
			16'h15b3: y = 16'h1ff;
			16'h15b4: y = 16'h1ff;
			16'h15b5: y = 16'h1ff;
			16'h15b6: y = 16'h1ff;
			16'h15b7: y = 16'h1ff;
			16'h15b8: y = 16'h1ff;
			16'h15b9: y = 16'h1ff;
			16'h15ba: y = 16'h1ff;
			16'h15bb: y = 16'h1ff;
			16'h15bc: y = 16'h1ff;
			16'h15bd: y = 16'h1ff;
			16'h15be: y = 16'h1ff;
			16'h15bf: y = 16'h1ff;
			16'h15c0: y = 16'h1ff;
			16'h15c1: y = 16'h1ff;
			16'h15c2: y = 16'h1ff;
			16'h15c3: y = 16'h1ff;
			16'h15c4: y = 16'h1ff;
			16'h15c5: y = 16'h1ff;
			16'h15c6: y = 16'h1ff;
			16'h15c7: y = 16'h1ff;
			16'h15c8: y = 16'h1ff;
			16'h15c9: y = 16'h1ff;
			16'h15ca: y = 16'h1ff;
			16'h15cb: y = 16'h1ff;
			16'h15cc: y = 16'h1ff;
			16'h15cd: y = 16'h1ff;
			16'h15ce: y = 16'h1ff;
			16'h15cf: y = 16'h1ff;
			16'h15d0: y = 16'h1ff;
			16'h15d1: y = 16'h1ff;
			16'h15d2: y = 16'h1ff;
			16'h15d3: y = 16'h1ff;
			16'h15d4: y = 16'h1ff;
			16'h15d5: y = 16'h1ff;
			16'h15d6: y = 16'h1ff;
			16'h15d7: y = 16'h1ff;
			16'h15d8: y = 16'h1ff;
			16'h15d9: y = 16'h1ff;
			16'h15da: y = 16'h1ff;
			16'h15db: y = 16'h1ff;
			16'h15dc: y = 16'h1ff;
			16'h15dd: y = 16'h1ff;
			16'h15de: y = 16'h1ff;
			16'h15df: y = 16'h1ff;
			16'h15e0: y = 16'h1ff;
			16'h15e1: y = 16'h1ff;
			16'h15e2: y = 16'h1ff;
			16'h15e3: y = 16'h1ff;
			16'h15e4: y = 16'h1ff;
			16'h15e5: y = 16'h1ff;
			16'h15e6: y = 16'h1ff;
			16'h15e7: y = 16'h1ff;
			16'h15e8: y = 16'h1ff;
			16'h15e9: y = 16'h1ff;
			16'h15ea: y = 16'h1ff;
			16'h15eb: y = 16'h1ff;
			16'h15ec: y = 16'h1ff;
			16'h15ed: y = 16'h1ff;
			16'h15ee: y = 16'h1ff;
			16'h15ef: y = 16'h1ff;
			16'h15f0: y = 16'h1ff;
			16'h15f1: y = 16'h1ff;
			16'h15f2: y = 16'h1ff;
			16'h15f3: y = 16'h1ff;
			16'h15f4: y = 16'h1ff;
			16'h15f5: y = 16'h1ff;
			16'h15f6: y = 16'h1ff;
			16'h15f7: y = 16'h1ff;
			16'h15f8: y = 16'h1ff;
			16'h15f9: y = 16'h1ff;
			16'h15fa: y = 16'h1ff;
			16'h15fb: y = 16'h1ff;
			16'h15fc: y = 16'h1ff;
			16'h15fd: y = 16'h1ff;
			16'h15fe: y = 16'h1ff;
			16'h15ff: y = 16'h1ff;
			16'h1600: y = 16'h1ff;
			16'h1601: y = 16'h1ff;
			16'h1602: y = 16'h1ff;
			16'h1603: y = 16'h1ff;
			16'h1604: y = 16'h1ff;
			16'h1605: y = 16'h1ff;
			16'h1606: y = 16'h1ff;
			16'h1607: y = 16'h1ff;
			16'h1608: y = 16'h1ff;
			16'h1609: y = 16'h1ff;
			16'h160a: y = 16'h1ff;
			16'h160b: y = 16'h1ff;
			16'h160c: y = 16'h1ff;
			16'h160d: y = 16'h1ff;
			16'h160e: y = 16'h1ff;
			16'h160f: y = 16'h1ff;
			16'h1610: y = 16'h1ff;
			16'h1611: y = 16'h1ff;
			16'h1612: y = 16'h1ff;
			16'h1613: y = 16'h1ff;
			16'h1614: y = 16'h1ff;
			16'h1615: y = 16'h1ff;
			16'h1616: y = 16'h1ff;
			16'h1617: y = 16'h1ff;
			16'h1618: y = 16'h1ff;
			16'h1619: y = 16'h1ff;
			16'h161a: y = 16'h1ff;
			16'h161b: y = 16'h1ff;
			16'h161c: y = 16'h1ff;
			16'h161d: y = 16'h1ff;
			16'h161e: y = 16'h1ff;
			16'h161f: y = 16'h1ff;
			16'h1620: y = 16'h1ff;
			16'h1621: y = 16'h1ff;
			16'h1622: y = 16'h1ff;
			16'h1623: y = 16'h1ff;
			16'h1624: y = 16'h1ff;
			16'h1625: y = 16'h1ff;
			16'h1626: y = 16'h1ff;
			16'h1627: y = 16'h1ff;
			16'h1628: y = 16'h1ff;
			16'h1629: y = 16'h1ff;
			16'h162a: y = 16'h1ff;
			16'h162b: y = 16'h1ff;
			16'h162c: y = 16'h1ff;
			16'h162d: y = 16'h1ff;
			16'h162e: y = 16'h1ff;
			16'h162f: y = 16'h1ff;
			16'h1630: y = 16'h1ff;
			16'h1631: y = 16'h1ff;
			16'h1632: y = 16'h1ff;
			16'h1633: y = 16'h1ff;
			16'h1634: y = 16'h1ff;
			16'h1635: y = 16'h1ff;
			16'h1636: y = 16'h1ff;
			16'h1637: y = 16'h1ff;
			16'h1638: y = 16'h1ff;
			16'h1639: y = 16'h1ff;
			16'h163a: y = 16'h1ff;
			16'h163b: y = 16'h1ff;
			16'h163c: y = 16'h1ff;
			16'h163d: y = 16'h1ff;
			16'h163e: y = 16'h1ff;
			16'h163f: y = 16'h1ff;
			16'h1640: y = 16'h1ff;
			16'h1641: y = 16'h1ff;
			16'h1642: y = 16'h1ff;
			16'h1643: y = 16'h1ff;
			16'h1644: y = 16'h1ff;
			16'h1645: y = 16'h1ff;
			16'h1646: y = 16'h1ff;
			16'h1647: y = 16'h1ff;
			16'h1648: y = 16'h1ff;
			16'h1649: y = 16'h1ff;
			16'h164a: y = 16'h1ff;
			16'h164b: y = 16'h1ff;
			16'h164c: y = 16'h1ff;
			16'h164d: y = 16'h1ff;
			16'h164e: y = 16'h1ff;
			16'h164f: y = 16'h1ff;
			16'h1650: y = 16'h1ff;
			16'h1651: y = 16'h1ff;
			16'h1652: y = 16'h1ff;
			16'h1653: y = 16'h1ff;
			16'h1654: y = 16'h1ff;
			16'h1655: y = 16'h1ff;
			16'h1656: y = 16'h1ff;
			16'h1657: y = 16'h1ff;
			16'h1658: y = 16'h1ff;
			16'h1659: y = 16'h1ff;
			16'h165a: y = 16'h1ff;
			16'h165b: y = 16'h1ff;
			16'h165c: y = 16'h1ff;
			16'h165d: y = 16'h1ff;
			16'h165e: y = 16'h1ff;
			16'h165f: y = 16'h1ff;
			16'h1660: y = 16'h1ff;
			16'h1661: y = 16'h1ff;
			16'h1662: y = 16'h1ff;
			16'h1663: y = 16'h1ff;
			16'h1664: y = 16'h1ff;
			16'h1665: y = 16'h1ff;
			16'h1666: y = 16'h1ff;
			16'h1667: y = 16'h1ff;
			16'h1668: y = 16'h1ff;
			16'h1669: y = 16'h1ff;
			16'h166a: y = 16'h1ff;
			16'h166b: y = 16'h1ff;
			16'h166c: y = 16'h1ff;
			16'h166d: y = 16'h1ff;
			16'h166e: y = 16'h1ff;
			16'h166f: y = 16'h1ff;
			16'h1670: y = 16'h1ff;
			16'h1671: y = 16'h1ff;
			16'h1672: y = 16'h1ff;
			16'h1673: y = 16'h1ff;
			16'h1674: y = 16'h1ff;
			16'h1675: y = 16'h1ff;
			16'h1676: y = 16'h1ff;
			16'h1677: y = 16'h1ff;
			16'h1678: y = 16'h1ff;
			16'h1679: y = 16'h1ff;
			16'h167a: y = 16'h1ff;
			16'h167b: y = 16'h1ff;
			16'h167c: y = 16'h1ff;
			16'h167d: y = 16'h1ff;
			16'h167e: y = 16'h1ff;
			16'h167f: y = 16'h1ff;
			16'h1680: y = 16'h1ff;
			16'h1681: y = 16'h1ff;
			16'h1682: y = 16'h1ff;
			16'h1683: y = 16'h1ff;
			16'h1684: y = 16'h1ff;
			16'h1685: y = 16'h1ff;
			16'h1686: y = 16'h1ff;
			16'h1687: y = 16'h1ff;
			16'h1688: y = 16'h1ff;
			16'h1689: y = 16'h1ff;
			16'h168a: y = 16'h1ff;
			16'h168b: y = 16'h1ff;
			16'h168c: y = 16'h1ff;
			16'h168d: y = 16'h1ff;
			16'h168e: y = 16'h1ff;
			16'h168f: y = 16'h1ff;
			16'h1690: y = 16'h1ff;
			16'h1691: y = 16'h1ff;
			16'h1692: y = 16'h1ff;
			16'h1693: y = 16'h1ff;
			16'h1694: y = 16'h1ff;
			16'h1695: y = 16'h1ff;
			16'h1696: y = 16'h1ff;
			16'h1697: y = 16'h1ff;
			16'h1698: y = 16'h1ff;
			16'h1699: y = 16'h1ff;
			16'h169a: y = 16'h1ff;
			16'h169b: y = 16'h1ff;
			16'h169c: y = 16'h1ff;
			16'h169d: y = 16'h1ff;
			16'h169e: y = 16'h1ff;
			16'h169f: y = 16'h1ff;
			16'h16a0: y = 16'h1ff;
			16'h16a1: y = 16'h1ff;
			16'h16a2: y = 16'h1ff;
			16'h16a3: y = 16'h1ff;
			16'h16a4: y = 16'h1ff;
			16'h16a5: y = 16'h1ff;
			16'h16a6: y = 16'h1ff;
			16'h16a7: y = 16'h1ff;
			16'h16a8: y = 16'h1ff;
			16'h16a9: y = 16'h1ff;
			16'h16aa: y = 16'h1ff;
			16'h16ab: y = 16'h1ff;
			16'h16ac: y = 16'h1ff;
			16'h16ad: y = 16'h1ff;
			16'h16ae: y = 16'h1ff;
			16'h16af: y = 16'h1ff;
			16'h16b0: y = 16'h1ff;
			16'h16b1: y = 16'h1ff;
			16'h16b2: y = 16'h1ff;
			16'h16b3: y = 16'h1ff;
			16'h16b4: y = 16'h1ff;
			16'h16b5: y = 16'h1ff;
			16'h16b6: y = 16'h1ff;
			16'h16b7: y = 16'h1ff;
			16'h16b8: y = 16'h1ff;
			16'h16b9: y = 16'h1ff;
			16'h16ba: y = 16'h1ff;
			16'h16bb: y = 16'h1ff;
			16'h16bc: y = 16'h1ff;
			16'h16bd: y = 16'h1ff;
			16'h16be: y = 16'h1ff;
			16'h16bf: y = 16'h1ff;
			16'h16c0: y = 16'h1ff;
			16'h16c1: y = 16'h1ff;
			16'h16c2: y = 16'h1ff;
			16'h16c3: y = 16'h1ff;
			16'h16c4: y = 16'h1ff;
			16'h16c5: y = 16'h1ff;
			16'h16c6: y = 16'h1ff;
			16'h16c7: y = 16'h1ff;
			16'h16c8: y = 16'h1ff;
			16'h16c9: y = 16'h1ff;
			16'h16ca: y = 16'h1ff;
			16'h16cb: y = 16'h1ff;
			16'h16cc: y = 16'h1ff;
			16'h16cd: y = 16'h1ff;
			16'h16ce: y = 16'h1ff;
			16'h16cf: y = 16'h1ff;
			16'h16d0: y = 16'h1ff;
			16'h16d1: y = 16'h1ff;
			16'h16d2: y = 16'h1ff;
			16'h16d3: y = 16'h1ff;
			16'h16d4: y = 16'h1ff;
			16'h16d5: y = 16'h1ff;
			16'h16d6: y = 16'h1ff;
			16'h16d7: y = 16'h1ff;
			16'h16d8: y = 16'h1ff;
			16'h16d9: y = 16'h1ff;
			16'h16da: y = 16'h1ff;
			16'h16db: y = 16'h1ff;
			16'h16dc: y = 16'h1ff;
			16'h16dd: y = 16'h1ff;
			16'h16de: y = 16'h1ff;
			16'h16df: y = 16'h1ff;
			16'h16e0: y = 16'h1ff;
			16'h16e1: y = 16'h1ff;
			16'h16e2: y = 16'h1ff;
			16'h16e3: y = 16'h1ff;
			16'h16e4: y = 16'h1ff;
			16'h16e5: y = 16'h1ff;
			16'h16e6: y = 16'h1ff;
			16'h16e7: y = 16'h1ff;
			16'h16e8: y = 16'h1ff;
			16'h16e9: y = 16'h1ff;
			16'h16ea: y = 16'h1ff;
			16'h16eb: y = 16'h1ff;
			16'h16ec: y = 16'h1ff;
			16'h16ed: y = 16'h1ff;
			16'h16ee: y = 16'h1ff;
			16'h16ef: y = 16'h1ff;
			16'h16f0: y = 16'h1ff;
			16'h16f1: y = 16'h1ff;
			16'h16f2: y = 16'h1ff;
			16'h16f3: y = 16'h1ff;
			16'h16f4: y = 16'h1ff;
			16'h16f5: y = 16'h1ff;
			16'h16f6: y = 16'h1ff;
			16'h16f7: y = 16'h1ff;
			16'h16f8: y = 16'h1ff;
			16'h16f9: y = 16'h1ff;
			16'h16fa: y = 16'h1ff;
			16'h16fb: y = 16'h1ff;
			16'h16fc: y = 16'h1ff;
			16'h16fd: y = 16'h1ff;
			16'h16fe: y = 16'h1ff;
			16'h16ff: y = 16'h1ff;
			16'h1700: y = 16'h1ff;
			16'h1701: y = 16'h1ff;
			16'h1702: y = 16'h1ff;
			16'h1703: y = 16'h1ff;
			16'h1704: y = 16'h1ff;
			16'h1705: y = 16'h1ff;
			16'h1706: y = 16'h1ff;
			16'h1707: y = 16'h1ff;
			16'h1708: y = 16'h1ff;
			16'h1709: y = 16'h1ff;
			16'h170a: y = 16'h1ff;
			16'h170b: y = 16'h1ff;
			16'h170c: y = 16'h1ff;
			16'h170d: y = 16'h1ff;
			16'h170e: y = 16'h1ff;
			16'h170f: y = 16'h1ff;
			16'h1710: y = 16'h1ff;
			16'h1711: y = 16'h1ff;
			16'h1712: y = 16'h1ff;
			16'h1713: y = 16'h1ff;
			16'h1714: y = 16'h1ff;
			16'h1715: y = 16'h1ff;
			16'h1716: y = 16'h1ff;
			16'h1717: y = 16'h1ff;
			16'h1718: y = 16'h1ff;
			16'h1719: y = 16'h1ff;
			16'h171a: y = 16'h1ff;
			16'h171b: y = 16'h1ff;
			16'h171c: y = 16'h1ff;
			16'h171d: y = 16'h1ff;
			16'h171e: y = 16'h1ff;
			16'h171f: y = 16'h1ff;
			16'h1720: y = 16'h1ff;
			16'h1721: y = 16'h1ff;
			16'h1722: y = 16'h1ff;
			16'h1723: y = 16'h1ff;
			16'h1724: y = 16'h1ff;
			16'h1725: y = 16'h1ff;
			16'h1726: y = 16'h1ff;
			16'h1727: y = 16'h1ff;
			16'h1728: y = 16'h1ff;
			16'h1729: y = 16'h1ff;
			16'h172a: y = 16'h1ff;
			16'h172b: y = 16'h1ff;
			16'h172c: y = 16'h1ff;
			16'h172d: y = 16'h1ff;
			16'h172e: y = 16'h1ff;
			16'h172f: y = 16'h1ff;
			16'h1730: y = 16'h1ff;
			16'h1731: y = 16'h1ff;
			16'h1732: y = 16'h1ff;
			16'h1733: y = 16'h1ff;
			16'h1734: y = 16'h1ff;
			16'h1735: y = 16'h1ff;
			16'h1736: y = 16'h1ff;
			16'h1737: y = 16'h1ff;
			16'h1738: y = 16'h1ff;
			16'h1739: y = 16'h1ff;
			16'h173a: y = 16'h1ff;
			16'h173b: y = 16'h1ff;
			16'h173c: y = 16'h1ff;
			16'h173d: y = 16'h1ff;
			16'h173e: y = 16'h1ff;
			16'h173f: y = 16'h1ff;
			16'h1740: y = 16'h1ff;
			16'h1741: y = 16'h1ff;
			16'h1742: y = 16'h1ff;
			16'h1743: y = 16'h1ff;
			16'h1744: y = 16'h1ff;
			16'h1745: y = 16'h1ff;
			16'h1746: y = 16'h1ff;
			16'h1747: y = 16'h1ff;
			16'h1748: y = 16'h1ff;
			16'h1749: y = 16'h1ff;
			16'h174a: y = 16'h1ff;
			16'h174b: y = 16'h1ff;
			16'h174c: y = 16'h1ff;
			16'h174d: y = 16'h1ff;
			16'h174e: y = 16'h1ff;
			16'h174f: y = 16'h1ff;
			16'h1750: y = 16'h1ff;
			16'h1751: y = 16'h1ff;
			16'h1752: y = 16'h1ff;
			16'h1753: y = 16'h1ff;
			16'h1754: y = 16'h1ff;
			16'h1755: y = 16'h1ff;
			16'h1756: y = 16'h1ff;
			16'h1757: y = 16'h1ff;
			16'h1758: y = 16'h1ff;
			16'h1759: y = 16'h1ff;
			16'h175a: y = 16'h1ff;
			16'h175b: y = 16'h1ff;
			16'h175c: y = 16'h1ff;
			16'h175d: y = 16'h1ff;
			16'h175e: y = 16'h1ff;
			16'h175f: y = 16'h1ff;
			16'h1760: y = 16'h1ff;
			16'h1761: y = 16'h1ff;
			16'h1762: y = 16'h1ff;
			16'h1763: y = 16'h1ff;
			16'h1764: y = 16'h1ff;
			16'h1765: y = 16'h1ff;
			16'h1766: y = 16'h1ff;
			16'h1767: y = 16'h1ff;
			16'h1768: y = 16'h1ff;
			16'h1769: y = 16'h1ff;
			16'h176a: y = 16'h1ff;
			16'h176b: y = 16'h1ff;
			16'h176c: y = 16'h1ff;
			16'h176d: y = 16'h1ff;
			16'h176e: y = 16'h1ff;
			16'h176f: y = 16'h1ff;
			16'h1770: y = 16'h1ff;
			16'h1771: y = 16'h1ff;
			16'h1772: y = 16'h1ff;
			16'h1773: y = 16'h1ff;
			16'h1774: y = 16'h1ff;
			16'h1775: y = 16'h1ff;
			16'h1776: y = 16'h1ff;
			16'h1777: y = 16'h1ff;
			16'h1778: y = 16'h1ff;
			16'h1779: y = 16'h1ff;
			16'h177a: y = 16'h1ff;
			16'h177b: y = 16'h1ff;
			16'h177c: y = 16'h1ff;
			16'h177d: y = 16'h1ff;
			16'h177e: y = 16'h1ff;
			16'h177f: y = 16'h1ff;
			16'h1780: y = 16'h1ff;
			16'h1781: y = 16'h1ff;
			16'h1782: y = 16'h1ff;
			16'h1783: y = 16'h1ff;
			16'h1784: y = 16'h1ff;
			16'h1785: y = 16'h1ff;
			16'h1786: y = 16'h1ff;
			16'h1787: y = 16'h1ff;
			16'h1788: y = 16'h1ff;
			16'h1789: y = 16'h1ff;
			16'h178a: y = 16'h1ff;
			16'h178b: y = 16'h1ff;
			16'h178c: y = 16'h1ff;
			16'h178d: y = 16'h1ff;
			16'h178e: y = 16'h1ff;
			16'h178f: y = 16'h1ff;
			16'h1790: y = 16'h1ff;
			16'h1791: y = 16'h1ff;
			16'h1792: y = 16'h1ff;
			16'h1793: y = 16'h1ff;
			16'h1794: y = 16'h1ff;
			16'h1795: y = 16'h1ff;
			16'h1796: y = 16'h1ff;
			16'h1797: y = 16'h1ff;
			16'h1798: y = 16'h1ff;
			16'h1799: y = 16'h1ff;
			16'h179a: y = 16'h1ff;
			16'h179b: y = 16'h1ff;
			16'h179c: y = 16'h1ff;
			16'h179d: y = 16'h1ff;
			16'h179e: y = 16'h1ff;
			16'h179f: y = 16'h1ff;
			16'h17a0: y = 16'h1ff;
			16'h17a1: y = 16'h1ff;
			16'h17a2: y = 16'h1ff;
			16'h17a3: y = 16'h1ff;
			16'h17a4: y = 16'h1ff;
			16'h17a5: y = 16'h1ff;
			16'h17a6: y = 16'h1ff;
			16'h17a7: y = 16'h1ff;
			16'h17a8: y = 16'h1ff;
			16'h17a9: y = 16'h1ff;
			16'h17aa: y = 16'h1ff;
			16'h17ab: y = 16'h1ff;
			16'h17ac: y = 16'h1ff;
			16'h17ad: y = 16'h1ff;
			16'h17ae: y = 16'h1ff;
			16'h17af: y = 16'h1ff;
			16'h17b0: y = 16'h1ff;
			16'h17b1: y = 16'h1ff;
			16'h17b2: y = 16'h1ff;
			16'h17b3: y = 16'h1ff;
			16'h17b4: y = 16'h1ff;
			16'h17b5: y = 16'h1ff;
			16'h17b6: y = 16'h1ff;
			16'h17b7: y = 16'h1ff;
			16'h17b8: y = 16'h1ff;
			16'h17b9: y = 16'h1ff;
			16'h17ba: y = 16'h1ff;
			16'h17bb: y = 16'h1ff;
			16'h17bc: y = 16'h1ff;
			16'h17bd: y = 16'h1ff;
			16'h17be: y = 16'h1ff;
			16'h17bf: y = 16'h1ff;
			16'h17c0: y = 16'h1ff;
			16'h17c1: y = 16'h1ff;
			16'h17c2: y = 16'h1ff;
			16'h17c3: y = 16'h1ff;
			16'h17c4: y = 16'h1ff;
			16'h17c5: y = 16'h1ff;
			16'h17c6: y = 16'h1ff;
			16'h17c7: y = 16'h1ff;
			16'h17c8: y = 16'h1ff;
			16'h17c9: y = 16'h1ff;
			16'h17ca: y = 16'h1ff;
			16'h17cb: y = 16'h1ff;
			16'h17cc: y = 16'h1ff;
			16'h17cd: y = 16'h1ff;
			16'h17ce: y = 16'h1ff;
			16'h17cf: y = 16'h1ff;
			16'h17d0: y = 16'h1ff;
			16'h17d1: y = 16'h1ff;
			16'h17d2: y = 16'h1ff;
			16'h17d3: y = 16'h1ff;
			16'h17d4: y = 16'h1ff;
			16'h17d5: y = 16'h1ff;
			16'h17d6: y = 16'h1ff;
			16'h17d7: y = 16'h1ff;
			16'h17d8: y = 16'h1ff;
			16'h17d9: y = 16'h1ff;
			16'h17da: y = 16'h1ff;
			16'h17db: y = 16'h1ff;
			16'h17dc: y = 16'h1ff;
			16'h17dd: y = 16'h1ff;
			16'h17de: y = 16'h1ff;
			16'h17df: y = 16'h1ff;
			16'h17e0: y = 16'h1ff;
			16'h17e1: y = 16'h1ff;
			16'h17e2: y = 16'h1ff;
			16'h17e3: y = 16'h1ff;
			16'h17e4: y = 16'h1ff;
			16'h17e5: y = 16'h1ff;
			16'h17e6: y = 16'h1ff;
			16'h17e7: y = 16'h1ff;
			16'h17e8: y = 16'h1ff;
			16'h17e9: y = 16'h1ff;
			16'h17ea: y = 16'h1ff;
			16'h17eb: y = 16'h1ff;
			16'h17ec: y = 16'h1ff;
			16'h17ed: y = 16'h1ff;
			16'h17ee: y = 16'h1ff;
			16'h17ef: y = 16'h1ff;
			16'h17f0: y = 16'h1ff;
			16'h17f1: y = 16'h1ff;
			16'h17f2: y = 16'h1ff;
			16'h17f3: y = 16'h1ff;
			16'h17f4: y = 16'h1ff;
			16'h17f5: y = 16'h1ff;
			16'h17f6: y = 16'h1ff;
			16'h17f7: y = 16'h1ff;
			16'h17f8: y = 16'h1ff;
			16'h17f9: y = 16'h1ff;
			16'h17fa: y = 16'h1ff;
			16'h17fb: y = 16'h1ff;
			16'h17fc: y = 16'h1ff;
			16'h17fd: y = 16'h1ff;
			16'h17fe: y = 16'h1ff;
			16'h17ff: y = 16'h1ff;
			16'h1800: y = 16'h1ff;
			16'h1801: y = 16'h1ff;
			16'h1802: y = 16'h1ff;
			16'h1803: y = 16'h1ff;
			16'h1804: y = 16'h1ff;
			16'h1805: y = 16'h1ff;
			16'h1806: y = 16'h1ff;
			16'h1807: y = 16'h1ff;
			16'h1808: y = 16'h1ff;
			16'h1809: y = 16'h1ff;
			16'h180a: y = 16'h1ff;
			16'h180b: y = 16'h1ff;
			16'h180c: y = 16'h1ff;
			16'h180d: y = 16'h1ff;
			16'h180e: y = 16'h1ff;
			16'h180f: y = 16'h1ff;
			16'h1810: y = 16'h1ff;
			16'h1811: y = 16'h1ff;
			16'h1812: y = 16'h1ff;
			16'h1813: y = 16'h1ff;
			16'h1814: y = 16'h1ff;
			16'h1815: y = 16'h1ff;
			16'h1816: y = 16'h1ff;
			16'h1817: y = 16'h1ff;
			16'h1818: y = 16'h1ff;
			16'h1819: y = 16'h1ff;
			16'h181a: y = 16'h1ff;
			16'h181b: y = 16'h1ff;
			16'h181c: y = 16'h1ff;
			16'h181d: y = 16'h1ff;
			16'h181e: y = 16'h1ff;
			16'h181f: y = 16'h1ff;
			16'h1820: y = 16'h1ff;
			16'h1821: y = 16'h1ff;
			16'h1822: y = 16'h1ff;
			16'h1823: y = 16'h1ff;
			16'h1824: y = 16'h1ff;
			16'h1825: y = 16'h1ff;
			16'h1826: y = 16'h1ff;
			16'h1827: y = 16'h1ff;
			16'h1828: y = 16'h1ff;
			16'h1829: y = 16'h1ff;
			16'h182a: y = 16'h1ff;
			16'h182b: y = 16'h1ff;
			16'h182c: y = 16'h1ff;
			16'h182d: y = 16'h1ff;
			16'h182e: y = 16'h1ff;
			16'h182f: y = 16'h1ff;
			16'h1830: y = 16'h1ff;
			16'h1831: y = 16'h1ff;
			16'h1832: y = 16'h1ff;
			16'h1833: y = 16'h1ff;
			16'h1834: y = 16'h1ff;
			16'h1835: y = 16'h1ff;
			16'h1836: y = 16'h1ff;
			16'h1837: y = 16'h1ff;
			16'h1838: y = 16'h1ff;
			16'h1839: y = 16'h1ff;
			16'h183a: y = 16'h1ff;
			16'h183b: y = 16'h1ff;
			16'h183c: y = 16'h1ff;
			16'h183d: y = 16'h1ff;
			16'h183e: y = 16'h1ff;
			16'h183f: y = 16'h1ff;
			16'h1840: y = 16'h1ff;
			16'h1841: y = 16'h1ff;
			16'h1842: y = 16'h1ff;
			16'h1843: y = 16'h1ff;
			16'h1844: y = 16'h1ff;
			16'h1845: y = 16'h1ff;
			16'h1846: y = 16'h1ff;
			16'h1847: y = 16'h1ff;
			16'h1848: y = 16'h1ff;
			16'h1849: y = 16'h1ff;
			16'h184a: y = 16'h1ff;
			16'h184b: y = 16'h1ff;
			16'h184c: y = 16'h1ff;
			16'h184d: y = 16'h1ff;
			16'h184e: y = 16'h1ff;
			16'h184f: y = 16'h1ff;
			16'h1850: y = 16'h1ff;
			16'h1851: y = 16'h1ff;
			16'h1852: y = 16'h1ff;
			16'h1853: y = 16'h1ff;
			16'h1854: y = 16'h1ff;
			16'h1855: y = 16'h1ff;
			16'h1856: y = 16'h1ff;
			16'h1857: y = 16'h1ff;
			16'h1858: y = 16'h1ff;
			16'h1859: y = 16'h1ff;
			16'h185a: y = 16'h1ff;
			16'h185b: y = 16'h1ff;
			16'h185c: y = 16'h1ff;
			16'h185d: y = 16'h1ff;
			16'h185e: y = 16'h1ff;
			16'h185f: y = 16'h1ff;
			16'h1860: y = 16'h1ff;
			16'h1861: y = 16'h1ff;
			16'h1862: y = 16'h1ff;
			16'h1863: y = 16'h1ff;
			16'h1864: y = 16'h1ff;
			16'h1865: y = 16'h1ff;
			16'h1866: y = 16'h1ff;
			16'h1867: y = 16'h1ff;
			16'h1868: y = 16'h1ff;
			16'h1869: y = 16'h1ff;
			16'h186a: y = 16'h1ff;
			16'h186b: y = 16'h1ff;
			16'h186c: y = 16'h1ff;
			16'h186d: y = 16'h1ff;
			16'h186e: y = 16'h1ff;
			16'h186f: y = 16'h1ff;
			16'h1870: y = 16'h1ff;
			16'h1871: y = 16'h1ff;
			16'h1872: y = 16'h1ff;
			16'h1873: y = 16'h1ff;
			16'h1874: y = 16'h1ff;
			16'h1875: y = 16'h1ff;
			16'h1876: y = 16'h1ff;
			16'h1877: y = 16'h1ff;
			16'h1878: y = 16'h1ff;
			16'h1879: y = 16'h1ff;
			16'h187a: y = 16'h1ff;
			16'h187b: y = 16'h1ff;
			16'h187c: y = 16'h1ff;
			16'h187d: y = 16'h1ff;
			16'h187e: y = 16'h1ff;
			16'h187f: y = 16'h1ff;
			16'h1880: y = 16'h1ff;
			16'h1881: y = 16'h1ff;
			16'h1882: y = 16'h1ff;
			16'h1883: y = 16'h1ff;
			16'h1884: y = 16'h1ff;
			16'h1885: y = 16'h1ff;
			16'h1886: y = 16'h1ff;
			16'h1887: y = 16'h1ff;
			16'h1888: y = 16'h1ff;
			16'h1889: y = 16'h1ff;
			16'h188a: y = 16'h1ff;
			16'h188b: y = 16'h1ff;
			16'h188c: y = 16'h1ff;
			16'h188d: y = 16'h1ff;
			16'h188e: y = 16'h1ff;
			16'h188f: y = 16'h1ff;
			16'h1890: y = 16'h1ff;
			16'h1891: y = 16'h1ff;
			16'h1892: y = 16'h1ff;
			16'h1893: y = 16'h1ff;
			16'h1894: y = 16'h1ff;
			16'h1895: y = 16'h1ff;
			16'h1896: y = 16'h1ff;
			16'h1897: y = 16'h1ff;
			16'h1898: y = 16'h1ff;
			16'h1899: y = 16'h1ff;
			16'h189a: y = 16'h1ff;
			16'h189b: y = 16'h1ff;
			16'h189c: y = 16'h1ff;
			16'h189d: y = 16'h1ff;
			16'h189e: y = 16'h1ff;
			16'h189f: y = 16'h1ff;
			16'h18a0: y = 16'h1ff;
			16'h18a1: y = 16'h1ff;
			16'h18a2: y = 16'h1ff;
			16'h18a3: y = 16'h1ff;
			16'h18a4: y = 16'h1ff;
			16'h18a5: y = 16'h1ff;
			16'h18a6: y = 16'h1ff;
			16'h18a7: y = 16'h1ff;
			16'h18a8: y = 16'h1ff;
			16'h18a9: y = 16'h1ff;
			16'h18aa: y = 16'h1ff;
			16'h18ab: y = 16'h1ff;
			16'h18ac: y = 16'h1ff;
			16'h18ad: y = 16'h1ff;
			16'h18ae: y = 16'h1ff;
			16'h18af: y = 16'h1ff;
			16'h18b0: y = 16'h1ff;
			16'h18b1: y = 16'h1ff;
			16'h18b2: y = 16'h1ff;
			16'h18b3: y = 16'h1ff;
			16'h18b4: y = 16'h1ff;
			16'h18b5: y = 16'h1ff;
			16'h18b6: y = 16'h1ff;
			16'h18b7: y = 16'h1ff;
			16'h18b8: y = 16'h1ff;
			16'h18b9: y = 16'h1ff;
			16'h18ba: y = 16'h1ff;
			16'h18bb: y = 16'h1ff;
			16'h18bc: y = 16'h1ff;
			16'h18bd: y = 16'h1ff;
			16'h18be: y = 16'h1ff;
			16'h18bf: y = 16'h1ff;
			16'h18c0: y = 16'h1ff;
			16'h18c1: y = 16'h1ff;
			16'h18c2: y = 16'h1ff;
			16'h18c3: y = 16'h1ff;
			16'h18c4: y = 16'h1ff;
			16'h18c5: y = 16'h1ff;
			16'h18c6: y = 16'h1ff;
			16'h18c7: y = 16'h1ff;
			16'h18c8: y = 16'h1ff;
			16'h18c9: y = 16'h1ff;
			16'h18ca: y = 16'h1ff;
			16'h18cb: y = 16'h1ff;
			16'h18cc: y = 16'h1ff;
			16'h18cd: y = 16'h1ff;
			16'h18ce: y = 16'h1ff;
			16'h18cf: y = 16'h1ff;
			16'h18d0: y = 16'h1ff;
			16'h18d1: y = 16'h1ff;
			16'h18d2: y = 16'h1ff;
			16'h18d3: y = 16'h1ff;
			16'h18d4: y = 16'h1ff;
			16'h18d5: y = 16'h1ff;
			16'h18d6: y = 16'h1ff;
			16'h18d7: y = 16'h1ff;
			16'h18d8: y = 16'h1ff;
			16'h18d9: y = 16'h1ff;
			16'h18da: y = 16'h1ff;
			16'h18db: y = 16'h1ff;
			16'h18dc: y = 16'h1ff;
			16'h18dd: y = 16'h1ff;
			16'h18de: y = 16'h1ff;
			16'h18df: y = 16'h1ff;
			16'h18e0: y = 16'h1ff;
			16'h18e1: y = 16'h1ff;
			16'h18e2: y = 16'h1ff;
			16'h18e3: y = 16'h1ff;
			16'h18e4: y = 16'h1ff;
			16'h18e5: y = 16'h1ff;
			16'h18e6: y = 16'h1ff;
			16'h18e7: y = 16'h1ff;
			16'h18e8: y = 16'h1ff;
			16'h18e9: y = 16'h1ff;
			16'h18ea: y = 16'h1ff;
			16'h18eb: y = 16'h1ff;
			16'h18ec: y = 16'h1ff;
			16'h18ed: y = 16'h1ff;
			16'h18ee: y = 16'h1ff;
			16'h18ef: y = 16'h1ff;
			16'h18f0: y = 16'h1ff;
			16'h18f1: y = 16'h1ff;
			16'h18f2: y = 16'h1ff;
			16'h18f3: y = 16'h1ff;
			16'h18f4: y = 16'h1ff;
			16'h18f5: y = 16'h1ff;
			16'h18f6: y = 16'h1ff;
			16'h18f7: y = 16'h1ff;
			16'h18f8: y = 16'h1ff;
			16'h18f9: y = 16'h1ff;
			16'h18fa: y = 16'h1ff;
			16'h18fb: y = 16'h1ff;
			16'h18fc: y = 16'h1ff;
			16'h18fd: y = 16'h1ff;
			16'h18fe: y = 16'h1ff;
			16'h18ff: y = 16'h1ff;
			16'h1900: y = 16'h1ff;
			16'h1901: y = 16'h1ff;
			16'h1902: y = 16'h1ff;
			16'h1903: y = 16'h1ff;
			16'h1904: y = 16'h1ff;
			16'h1905: y = 16'h1ff;
			16'h1906: y = 16'h1ff;
			16'h1907: y = 16'h1ff;
			16'h1908: y = 16'h1ff;
			16'h1909: y = 16'h1ff;
			16'h190a: y = 16'h1ff;
			16'h190b: y = 16'h1ff;
			16'h190c: y = 16'h1ff;
			16'h190d: y = 16'h1ff;
			16'h190e: y = 16'h1ff;
			16'h190f: y = 16'h1ff;
			16'h1910: y = 16'h1ff;
			16'h1911: y = 16'h1ff;
			16'h1912: y = 16'h1ff;
			16'h1913: y = 16'h1ff;
			16'h1914: y = 16'h1ff;
			16'h1915: y = 16'h1ff;
			16'h1916: y = 16'h1ff;
			16'h1917: y = 16'h1ff;
			16'h1918: y = 16'h1ff;
			16'h1919: y = 16'h1ff;
			16'h191a: y = 16'h1ff;
			16'h191b: y = 16'h1ff;
			16'h191c: y = 16'h1ff;
			16'h191d: y = 16'h1ff;
			16'h191e: y = 16'h1ff;
			16'h191f: y = 16'h1ff;
			16'h1920: y = 16'h1ff;
			16'h1921: y = 16'h1ff;
			16'h1922: y = 16'h1ff;
			16'h1923: y = 16'h1ff;
			16'h1924: y = 16'h1ff;
			16'h1925: y = 16'h1ff;
			16'h1926: y = 16'h1ff;
			16'h1927: y = 16'h1ff;
			16'h1928: y = 16'h1ff;
			16'h1929: y = 16'h1ff;
			16'h192a: y = 16'h1ff;
			16'h192b: y = 16'h1ff;
			16'h192c: y = 16'h1ff;
			16'h192d: y = 16'h1ff;
			16'h192e: y = 16'h1ff;
			16'h192f: y = 16'h1ff;
			16'h1930: y = 16'h1ff;
			16'h1931: y = 16'h1ff;
			16'h1932: y = 16'h1ff;
			16'h1933: y = 16'h1ff;
			16'h1934: y = 16'h1ff;
			16'h1935: y = 16'h1ff;
			16'h1936: y = 16'h1ff;
			16'h1937: y = 16'h1ff;
			16'h1938: y = 16'h1ff;
			16'h1939: y = 16'h1ff;
			16'h193a: y = 16'h1ff;
			16'h193b: y = 16'h1ff;
			16'h193c: y = 16'h1ff;
			16'h193d: y = 16'h1ff;
			16'h193e: y = 16'h1ff;
			16'h193f: y = 16'h1ff;
			16'h1940: y = 16'h1ff;
			16'h1941: y = 16'h1ff;
			16'h1942: y = 16'h1ff;
			16'h1943: y = 16'h1ff;
			16'h1944: y = 16'h1ff;
			16'h1945: y = 16'h1ff;
			16'h1946: y = 16'h1ff;
			16'h1947: y = 16'h1ff;
			16'h1948: y = 16'h1ff;
			16'h1949: y = 16'h1ff;
			16'h194a: y = 16'h1ff;
			16'h194b: y = 16'h1ff;
			16'h194c: y = 16'h1ff;
			16'h194d: y = 16'h1ff;
			16'h194e: y = 16'h1ff;
			16'h194f: y = 16'h1ff;
			16'h1950: y = 16'h1ff;
			16'h1951: y = 16'h1ff;
			16'h1952: y = 16'h1ff;
			16'h1953: y = 16'h1ff;
			16'h1954: y = 16'h1ff;
			16'h1955: y = 16'h1ff;
			16'h1956: y = 16'h1ff;
			16'h1957: y = 16'h1ff;
			16'h1958: y = 16'h1ff;
			16'h1959: y = 16'h1ff;
			16'h195a: y = 16'h1ff;
			16'h195b: y = 16'h1ff;
			16'h195c: y = 16'h1ff;
			16'h195d: y = 16'h1ff;
			16'h195e: y = 16'h1ff;
			16'h195f: y = 16'h1ff;
			16'h1960: y = 16'h1ff;
			16'h1961: y = 16'h1ff;
			16'h1962: y = 16'h1ff;
			16'h1963: y = 16'h1ff;
			16'h1964: y = 16'h1ff;
			16'h1965: y = 16'h1ff;
			16'h1966: y = 16'h1ff;
			16'h1967: y = 16'h1ff;
			16'h1968: y = 16'h1ff;
			16'h1969: y = 16'h1ff;
			16'h196a: y = 16'h1ff;
			16'h196b: y = 16'h1ff;
			16'h196c: y = 16'h1ff;
			16'h196d: y = 16'h1ff;
			16'h196e: y = 16'h1ff;
			16'h196f: y = 16'h1ff;
			16'h1970: y = 16'h1ff;
			16'h1971: y = 16'h1ff;
			16'h1972: y = 16'h1ff;
			16'h1973: y = 16'h1ff;
			16'h1974: y = 16'h1ff;
			16'h1975: y = 16'h1ff;
			16'h1976: y = 16'h1ff;
			16'h1977: y = 16'h1ff;
			16'h1978: y = 16'h1ff;
			16'h1979: y = 16'h1ff;
			16'h197a: y = 16'h1ff;
			16'h197b: y = 16'h1ff;
			16'h197c: y = 16'h1ff;
			16'h197d: y = 16'h1ff;
			16'h197e: y = 16'h1ff;
			16'h197f: y = 16'h1ff;
			16'h1980: y = 16'h1ff;
			16'h1981: y = 16'h1ff;
			16'h1982: y = 16'h1ff;
			16'h1983: y = 16'h1ff;
			16'h1984: y = 16'h1ff;
			16'h1985: y = 16'h1ff;
			16'h1986: y = 16'h1ff;
			16'h1987: y = 16'h1ff;
			16'h1988: y = 16'h1ff;
			16'h1989: y = 16'h1ff;
			16'h198a: y = 16'h1ff;
			16'h198b: y = 16'h1ff;
			16'h198c: y = 16'h1ff;
			16'h198d: y = 16'h1ff;
			16'h198e: y = 16'h1ff;
			16'h198f: y = 16'h1ff;
			16'h1990: y = 16'h1ff;
			16'h1991: y = 16'h1ff;
			16'h1992: y = 16'h1ff;
			16'h1993: y = 16'h1ff;
			16'h1994: y = 16'h1ff;
			16'h1995: y = 16'h1ff;
			16'h1996: y = 16'h1ff;
			16'h1997: y = 16'h1ff;
			16'h1998: y = 16'h1ff;
			16'h1999: y = 16'h1ff;
			16'h199a: y = 16'h1ff;
			16'h199b: y = 16'h1ff;
			16'h199c: y = 16'h1ff;
			16'h199d: y = 16'h1ff;
			16'h199e: y = 16'h1ff;
			16'h199f: y = 16'h1ff;
			16'h19a0: y = 16'h1ff;
			16'h19a1: y = 16'h1ff;
			16'h19a2: y = 16'h1ff;
			16'h19a3: y = 16'h1ff;
			16'h19a4: y = 16'h1ff;
			16'h19a5: y = 16'h1ff;
			16'h19a6: y = 16'h1ff;
			16'h19a7: y = 16'h1ff;
			16'h19a8: y = 16'h1ff;
			16'h19a9: y = 16'h1ff;
			16'h19aa: y = 16'h1ff;
			16'h19ab: y = 16'h1ff;
			16'h19ac: y = 16'h1ff;
			16'h19ad: y = 16'h1ff;
			16'h19ae: y = 16'h1ff;
			16'h19af: y = 16'h1ff;
			16'h19b0: y = 16'h1ff;
			16'h19b1: y = 16'h1ff;
			16'h19b2: y = 16'h1ff;
			16'h19b3: y = 16'h1ff;
			16'h19b4: y = 16'h1ff;
			16'h19b5: y = 16'h1ff;
			16'h19b6: y = 16'h1ff;
			16'h19b7: y = 16'h1ff;
			16'h19b8: y = 16'h1ff;
			16'h19b9: y = 16'h1ff;
			16'h19ba: y = 16'h1ff;
			16'h19bb: y = 16'h1ff;
			16'h19bc: y = 16'h1ff;
			16'h19bd: y = 16'h1ff;
			16'h19be: y = 16'h1ff;
			16'h19bf: y = 16'h1ff;
			16'h19c0: y = 16'h1ff;
			16'h19c1: y = 16'h1ff;
			16'h19c2: y = 16'h1ff;
			16'h19c3: y = 16'h1ff;
			16'h19c4: y = 16'h1ff;
			16'h19c5: y = 16'h1ff;
			16'h19c6: y = 16'h1ff;
			16'h19c7: y = 16'h1ff;
			16'h19c8: y = 16'h1ff;
			16'h19c9: y = 16'h1ff;
			16'h19ca: y = 16'h1ff;
			16'h19cb: y = 16'h1ff;
			16'h19cc: y = 16'h1ff;
			16'h19cd: y = 16'h1ff;
			16'h19ce: y = 16'h1ff;
			16'h19cf: y = 16'h1ff;
			16'h19d0: y = 16'h1ff;
			16'h19d1: y = 16'h1ff;
			16'h19d2: y = 16'h1ff;
			16'h19d3: y = 16'h1ff;
			16'h19d4: y = 16'h1ff;
			16'h19d5: y = 16'h1ff;
			16'h19d6: y = 16'h1ff;
			16'h19d7: y = 16'h1ff;
			16'h19d8: y = 16'h1ff;
			16'h19d9: y = 16'h1ff;
			16'h19da: y = 16'h1ff;
			16'h19db: y = 16'h1ff;
			16'h19dc: y = 16'h1ff;
			16'h19dd: y = 16'h1ff;
			16'h19de: y = 16'h1ff;
			16'h19df: y = 16'h1ff;
			16'h19e0: y = 16'h1ff;
			16'h19e1: y = 16'h1ff;
			16'h19e2: y = 16'h1ff;
			16'h19e3: y = 16'h1ff;
			16'h19e4: y = 16'h1ff;
			16'h19e5: y = 16'h1ff;
			16'h19e6: y = 16'h1ff;
			16'h19e7: y = 16'h1ff;
			16'h19e8: y = 16'h1ff;
			16'h19e9: y = 16'h1ff;
			16'h19ea: y = 16'h1ff;
			16'h19eb: y = 16'h1ff;
			16'h19ec: y = 16'h1ff;
			16'h19ed: y = 16'h1ff;
			16'h19ee: y = 16'h1ff;
			16'h19ef: y = 16'h1ff;
			16'h19f0: y = 16'h1ff;
			16'h19f1: y = 16'h1ff;
			16'h19f2: y = 16'h1ff;
			16'h19f3: y = 16'h1ff;
			16'h19f4: y = 16'h1ff;
			16'h19f5: y = 16'h1ff;
			16'h19f6: y = 16'h1ff;
			16'h19f7: y = 16'h1ff;
			16'h19f8: y = 16'h1ff;
			16'h19f9: y = 16'h1ff;
			16'h19fa: y = 16'h1ff;
			16'h19fb: y = 16'h1ff;
			16'h19fc: y = 16'h1ff;
			16'h19fd: y = 16'h1ff;
			16'h19fe: y = 16'h1ff;
			16'h19ff: y = 16'h1ff;
			16'h1a00: y = 16'h1ff;
			16'h1a01: y = 16'h1ff;
			16'h1a02: y = 16'h1ff;
			16'h1a03: y = 16'h1ff;
			16'h1a04: y = 16'h1ff;
			16'h1a05: y = 16'h1ff;
			16'h1a06: y = 16'h1ff;
			16'h1a07: y = 16'h1ff;
			16'h1a08: y = 16'h1ff;
			16'h1a09: y = 16'h1ff;
			16'h1a0a: y = 16'h1ff;
			16'h1a0b: y = 16'h1ff;
			16'h1a0c: y = 16'h1ff;
			16'h1a0d: y = 16'h1ff;
			16'h1a0e: y = 16'h1ff;
			16'h1a0f: y = 16'h1ff;
			16'h1a10: y = 16'h1ff;
			16'h1a11: y = 16'h1ff;
			16'h1a12: y = 16'h1ff;
			16'h1a13: y = 16'h1ff;
			16'h1a14: y = 16'h1ff;
			16'h1a15: y = 16'h1ff;
			16'h1a16: y = 16'h1ff;
			16'h1a17: y = 16'h1ff;
			16'h1a18: y = 16'h1ff;
			16'h1a19: y = 16'h1ff;
			16'h1a1a: y = 16'h1ff;
			16'h1a1b: y = 16'h1ff;
			16'h1a1c: y = 16'h1ff;
			16'h1a1d: y = 16'h1ff;
			16'h1a1e: y = 16'h1ff;
			16'h1a1f: y = 16'h1ff;
			16'h1a20: y = 16'h1ff;
			16'h1a21: y = 16'h1ff;
			16'h1a22: y = 16'h1ff;
			16'h1a23: y = 16'h1ff;
			16'h1a24: y = 16'h1ff;
			16'h1a25: y = 16'h1ff;
			16'h1a26: y = 16'h1ff;
			16'h1a27: y = 16'h1ff;
			16'h1a28: y = 16'h1ff;
			16'h1a29: y = 16'h1ff;
			16'h1a2a: y = 16'h1ff;
			16'h1a2b: y = 16'h1ff;
			16'h1a2c: y = 16'h1ff;
			16'h1a2d: y = 16'h1ff;
			16'h1a2e: y = 16'h1ff;
			16'h1a2f: y = 16'h1ff;
			16'h1a30: y = 16'h1ff;
			16'h1a31: y = 16'h1ff;
			16'h1a32: y = 16'h1ff;
			16'h1a33: y = 16'h1ff;
			16'h1a34: y = 16'h1ff;
			16'h1a35: y = 16'h1ff;
			16'h1a36: y = 16'h1ff;
			16'h1a37: y = 16'h1ff;
			16'h1a38: y = 16'h1ff;
			16'h1a39: y = 16'h1ff;
			16'h1a3a: y = 16'h1ff;
			16'h1a3b: y = 16'h1ff;
			16'h1a3c: y = 16'h1ff;
			16'h1a3d: y = 16'h1ff;
			16'h1a3e: y = 16'h1ff;
			16'h1a3f: y = 16'h1ff;
			16'h1a40: y = 16'h1ff;
			16'h1a41: y = 16'h1ff;
			16'h1a42: y = 16'h1ff;
			16'h1a43: y = 16'h1ff;
			16'h1a44: y = 16'h1ff;
			16'h1a45: y = 16'h1ff;
			16'h1a46: y = 16'h1ff;
			16'h1a47: y = 16'h1ff;
			16'h1a48: y = 16'h1ff;
			16'h1a49: y = 16'h1ff;
			16'h1a4a: y = 16'h1ff;
			16'h1a4b: y = 16'h1ff;
			16'h1a4c: y = 16'h1ff;
			16'h1a4d: y = 16'h1ff;
			16'h1a4e: y = 16'h1ff;
			16'h1a4f: y = 16'h1ff;
			16'h1a50: y = 16'h1ff;
			16'h1a51: y = 16'h1ff;
			16'h1a52: y = 16'h1ff;
			16'h1a53: y = 16'h1ff;
			16'h1a54: y = 16'h1ff;
			16'h1a55: y = 16'h1ff;
			16'h1a56: y = 16'h1ff;
			16'h1a57: y = 16'h1ff;
			16'h1a58: y = 16'h1ff;
			16'h1a59: y = 16'h1ff;
			16'h1a5a: y = 16'h1ff;
			16'h1a5b: y = 16'h1ff;
			16'h1a5c: y = 16'h1ff;
			16'h1a5d: y = 16'h1ff;
			16'h1a5e: y = 16'h1ff;
			16'h1a5f: y = 16'h1ff;
			16'h1a60: y = 16'h1ff;
			16'h1a61: y = 16'h1ff;
			16'h1a62: y = 16'h1ff;
			16'h1a63: y = 16'h1ff;
			16'h1a64: y = 16'h1ff;
			16'h1a65: y = 16'h1ff;
			16'h1a66: y = 16'h1ff;
			16'h1a67: y = 16'h1ff;
			16'h1a68: y = 16'h1ff;
			16'h1a69: y = 16'h1ff;
			16'h1a6a: y = 16'h1ff;
			16'h1a6b: y = 16'h1ff;
			16'h1a6c: y = 16'h1ff;
			16'h1a6d: y = 16'h1ff;
			16'h1a6e: y = 16'h1ff;
			16'h1a6f: y = 16'h1ff;
			16'h1a70: y = 16'h1ff;
			16'h1a71: y = 16'h1ff;
			16'h1a72: y = 16'h1ff;
			16'h1a73: y = 16'h1ff;
			16'h1a74: y = 16'h1ff;
			16'h1a75: y = 16'h1ff;
			16'h1a76: y = 16'h1ff;
			16'h1a77: y = 16'h1ff;
			16'h1a78: y = 16'h1ff;
			16'h1a79: y = 16'h1ff;
			16'h1a7a: y = 16'h1ff;
			16'h1a7b: y = 16'h1ff;
			16'h1a7c: y = 16'h1ff;
			16'h1a7d: y = 16'h1ff;
			16'h1a7e: y = 16'h1ff;
			16'h1a7f: y = 16'h1ff;
			16'h1a80: y = 16'h1ff;
			16'h1a81: y = 16'h1ff;
			16'h1a82: y = 16'h1ff;
			16'h1a83: y = 16'h1ff;
			16'h1a84: y = 16'h1ff;
			16'h1a85: y = 16'h1ff;
			16'h1a86: y = 16'h1ff;
			16'h1a87: y = 16'h1ff;
			16'h1a88: y = 16'h1ff;
			16'h1a89: y = 16'h1ff;
			16'h1a8a: y = 16'h1ff;
			16'h1a8b: y = 16'h1ff;
			16'h1a8c: y = 16'h1ff;
			16'h1a8d: y = 16'h1ff;
			16'h1a8e: y = 16'h1ff;
			16'h1a8f: y = 16'h1ff;
			16'h1a90: y = 16'h1ff;
			16'h1a91: y = 16'h1ff;
			16'h1a92: y = 16'h1ff;
			16'h1a93: y = 16'h1ff;
			16'h1a94: y = 16'h1ff;
			16'h1a95: y = 16'h1ff;
			16'h1a96: y = 16'h1ff;
			16'h1a97: y = 16'h1ff;
			16'h1a98: y = 16'h1ff;
			16'h1a99: y = 16'h1ff;
			16'h1a9a: y = 16'h1ff;
			16'h1a9b: y = 16'h1ff;
			16'h1a9c: y = 16'h1ff;
			16'h1a9d: y = 16'h1ff;
			16'h1a9e: y = 16'h1ff;
			16'h1a9f: y = 16'h1ff;
			16'h1aa0: y = 16'h1ff;
			16'h1aa1: y = 16'h1ff;
			16'h1aa2: y = 16'h1ff;
			16'h1aa3: y = 16'h1ff;
			16'h1aa4: y = 16'h1ff;
			16'h1aa5: y = 16'h1ff;
			16'h1aa6: y = 16'h1ff;
			16'h1aa7: y = 16'h1ff;
			16'h1aa8: y = 16'h1ff;
			16'h1aa9: y = 16'h1ff;
			16'h1aaa: y = 16'h1ff;
			16'h1aab: y = 16'h1ff;
			16'h1aac: y = 16'h1ff;
			16'h1aad: y = 16'h1ff;
			16'h1aae: y = 16'h1ff;
			16'h1aaf: y = 16'h1ff;
			16'h1ab0: y = 16'h1ff;
			16'h1ab1: y = 16'h1ff;
			16'h1ab2: y = 16'h1ff;
			16'h1ab3: y = 16'h1ff;
			16'h1ab4: y = 16'h1ff;
			16'h1ab5: y = 16'h1ff;
			16'h1ab6: y = 16'h1ff;
			16'h1ab7: y = 16'h1ff;
			16'h1ab8: y = 16'h1ff;
			16'h1ab9: y = 16'h1ff;
			16'h1aba: y = 16'h1ff;
			16'h1abb: y = 16'h1ff;
			16'h1abc: y = 16'h1ff;
			16'h1abd: y = 16'h1ff;
			16'h1abe: y = 16'h1ff;
			16'h1abf: y = 16'h1ff;
			16'h1ac0: y = 16'h1ff;
			16'h1ac1: y = 16'h1ff;
			16'h1ac2: y = 16'h1ff;
			16'h1ac3: y = 16'h1ff;
			16'h1ac4: y = 16'h1ff;
			16'h1ac5: y = 16'h1ff;
			16'h1ac6: y = 16'h1ff;
			16'h1ac7: y = 16'h1ff;
			16'h1ac8: y = 16'h1ff;
			16'h1ac9: y = 16'h1ff;
			16'h1aca: y = 16'h1ff;
			16'h1acb: y = 16'h1ff;
			16'h1acc: y = 16'h1ff;
			16'h1acd: y = 16'h1ff;
			16'h1ace: y = 16'h1ff;
			16'h1acf: y = 16'h1ff;
			16'h1ad0: y = 16'h1ff;
			16'h1ad1: y = 16'h1ff;
			16'h1ad2: y = 16'h1ff;
			16'h1ad3: y = 16'h1ff;
			16'h1ad4: y = 16'h1ff;
			16'h1ad5: y = 16'h1ff;
			16'h1ad6: y = 16'h1ff;
			16'h1ad7: y = 16'h1ff;
			16'h1ad8: y = 16'h1ff;
			16'h1ad9: y = 16'h1ff;
			16'h1ada: y = 16'h1ff;
			16'h1adb: y = 16'h1ff;
			16'h1adc: y = 16'h1ff;
			16'h1add: y = 16'h1ff;
			16'h1ade: y = 16'h1ff;
			16'h1adf: y = 16'h1ff;
			16'h1ae0: y = 16'h1ff;
			16'h1ae1: y = 16'h1ff;
			16'h1ae2: y = 16'h1ff;
			16'h1ae3: y = 16'h1ff;
			16'h1ae4: y = 16'h1ff;
			16'h1ae5: y = 16'h1ff;
			16'h1ae6: y = 16'h1ff;
			16'h1ae7: y = 16'h1ff;
			16'h1ae8: y = 16'h1ff;
			16'h1ae9: y = 16'h1ff;
			16'h1aea: y = 16'h1ff;
			16'h1aeb: y = 16'h1ff;
			16'h1aec: y = 16'h1ff;
			16'h1aed: y = 16'h1ff;
			16'h1aee: y = 16'h1ff;
			16'h1aef: y = 16'h1ff;
			16'h1af0: y = 16'h1ff;
			16'h1af1: y = 16'h1ff;
			16'h1af2: y = 16'h1ff;
			16'h1af3: y = 16'h1ff;
			16'h1af4: y = 16'h1ff;
			16'h1af5: y = 16'h1ff;
			16'h1af6: y = 16'h1ff;
			16'h1af7: y = 16'h1ff;
			16'h1af8: y = 16'h1ff;
			16'h1af9: y = 16'h1ff;
			16'h1afa: y = 16'h1ff;
			16'h1afb: y = 16'h1ff;
			16'h1afc: y = 16'h1ff;
			16'h1afd: y = 16'h1ff;
			16'h1afe: y = 16'h1ff;
			16'h1aff: y = 16'h1ff;
			16'h1b00: y = 16'h1ff;
			16'h1b01: y = 16'h1ff;
			16'h1b02: y = 16'h1ff;
			16'h1b03: y = 16'h1ff;
			16'h1b04: y = 16'h1ff;
			16'h1b05: y = 16'h1ff;
			16'h1b06: y = 16'h1ff;
			16'h1b07: y = 16'h1ff;
			16'h1b08: y = 16'h1ff;
			16'h1b09: y = 16'h1ff;
			16'h1b0a: y = 16'h1ff;
			16'h1b0b: y = 16'h1ff;
			16'h1b0c: y = 16'h1ff;
			16'h1b0d: y = 16'h1ff;
			16'h1b0e: y = 16'h1ff;
			16'h1b0f: y = 16'h1ff;
			16'h1b10: y = 16'h1ff;
			16'h1b11: y = 16'h1ff;
			16'h1b12: y = 16'h1ff;
			16'h1b13: y = 16'h1ff;
			16'h1b14: y = 16'h1ff;
			16'h1b15: y = 16'h1ff;
			16'h1b16: y = 16'h1ff;
			16'h1b17: y = 16'h1ff;
			16'h1b18: y = 16'h1ff;
			16'h1b19: y = 16'h1ff;
			16'h1b1a: y = 16'h1ff;
			16'h1b1b: y = 16'h1ff;
			16'h1b1c: y = 16'h1ff;
			16'h1b1d: y = 16'h1ff;
			16'h1b1e: y = 16'h1ff;
			16'h1b1f: y = 16'h1ff;
			16'h1b20: y = 16'h1ff;
			16'h1b21: y = 16'h1ff;
			16'h1b22: y = 16'h1ff;
			16'h1b23: y = 16'h1ff;
			16'h1b24: y = 16'h1ff;
			16'h1b25: y = 16'h1ff;
			16'h1b26: y = 16'h1ff;
			16'h1b27: y = 16'h1ff;
			16'h1b28: y = 16'h1ff;
			16'h1b29: y = 16'h1ff;
			16'h1b2a: y = 16'h1ff;
			16'h1b2b: y = 16'h1ff;
			16'h1b2c: y = 16'h1ff;
			16'h1b2d: y = 16'h1ff;
			16'h1b2e: y = 16'h1ff;
			16'h1b2f: y = 16'h1ff;
			16'h1b30: y = 16'h1ff;
			16'h1b31: y = 16'h1ff;
			16'h1b32: y = 16'h1ff;
			16'h1b33: y = 16'h1ff;
			16'h1b34: y = 16'h1ff;
			16'h1b35: y = 16'h1ff;
			16'h1b36: y = 16'h1ff;
			16'h1b37: y = 16'h1ff;
			16'h1b38: y = 16'h1ff;
			16'h1b39: y = 16'h1ff;
			16'h1b3a: y = 16'h1ff;
			16'h1b3b: y = 16'h1ff;
			16'h1b3c: y = 16'h1ff;
			16'h1b3d: y = 16'h1ff;
			16'h1b3e: y = 16'h1ff;
			16'h1b3f: y = 16'h1ff;
			16'h1b40: y = 16'h1ff;
			16'h1b41: y = 16'h1ff;
			16'h1b42: y = 16'h1ff;
			16'h1b43: y = 16'h1ff;
			16'h1b44: y = 16'h1ff;
			16'h1b45: y = 16'h1ff;
			16'h1b46: y = 16'h1ff;
			16'h1b47: y = 16'h1ff;
			16'h1b48: y = 16'h1ff;
			16'h1b49: y = 16'h1ff;
			16'h1b4a: y = 16'h1ff;
			16'h1b4b: y = 16'h1ff;
			16'h1b4c: y = 16'h1ff;
			16'h1b4d: y = 16'h1ff;
			16'h1b4e: y = 16'h1ff;
			16'h1b4f: y = 16'h1ff;
			16'h1b50: y = 16'h1ff;
			16'h1b51: y = 16'h1ff;
			16'h1b52: y = 16'h1ff;
			16'h1b53: y = 16'h1ff;
			16'h1b54: y = 16'h1ff;
			16'h1b55: y = 16'h1ff;
			16'h1b56: y = 16'h1ff;
			16'h1b57: y = 16'h1ff;
			16'h1b58: y = 16'h1ff;
			16'h1b59: y = 16'h1ff;
			16'h1b5a: y = 16'h1ff;
			16'h1b5b: y = 16'h1ff;
			16'h1b5c: y = 16'h1ff;
			16'h1b5d: y = 16'h1ff;
			16'h1b5e: y = 16'h1ff;
			16'h1b5f: y = 16'h1ff;
			16'h1b60: y = 16'h1ff;
			16'h1b61: y = 16'h1ff;
			16'h1b62: y = 16'h1ff;
			16'h1b63: y = 16'h1ff;
			16'h1b64: y = 16'h1ff;
			16'h1b65: y = 16'h1ff;
			16'h1b66: y = 16'h1ff;
			16'h1b67: y = 16'h1ff;
			16'h1b68: y = 16'h1ff;
			16'h1b69: y = 16'h1ff;
			16'h1b6a: y = 16'h1ff;
			16'h1b6b: y = 16'h1ff;
			16'h1b6c: y = 16'h1ff;
			16'h1b6d: y = 16'h1ff;
			16'h1b6e: y = 16'h1ff;
			16'h1b6f: y = 16'h1ff;
			16'h1b70: y = 16'h1ff;
			16'h1b71: y = 16'h1ff;
			16'h1b72: y = 16'h1ff;
			16'h1b73: y = 16'h1ff;
			16'h1b74: y = 16'h1ff;
			16'h1b75: y = 16'h1ff;
			16'h1b76: y = 16'h1ff;
			16'h1b77: y = 16'h1ff;
			16'h1b78: y = 16'h1ff;
			16'h1b79: y = 16'h1ff;
			16'h1b7a: y = 16'h1ff;
			16'h1b7b: y = 16'h1ff;
			16'h1b7c: y = 16'h1ff;
			16'h1b7d: y = 16'h1ff;
			16'h1b7e: y = 16'h1ff;
			16'h1b7f: y = 16'h1ff;
			16'h1b80: y = 16'h1ff;
			16'h1b81: y = 16'h1ff;
			16'h1b82: y = 16'h1ff;
			16'h1b83: y = 16'h1ff;
			16'h1b84: y = 16'h1ff;
			16'h1b85: y = 16'h1ff;
			16'h1b86: y = 16'h1ff;
			16'h1b87: y = 16'h1ff;
			16'h1b88: y = 16'h1ff;
			16'h1b89: y = 16'h1ff;
			16'h1b8a: y = 16'h1ff;
			16'h1b8b: y = 16'h1ff;
			16'h1b8c: y = 16'h1ff;
			16'h1b8d: y = 16'h1ff;
			16'h1b8e: y = 16'h1ff;
			16'h1b8f: y = 16'h1ff;
			16'h1b90: y = 16'h1ff;
			16'h1b91: y = 16'h1ff;
			16'h1b92: y = 16'h1ff;
			16'h1b93: y = 16'h1ff;
			16'h1b94: y = 16'h1ff;
			16'h1b95: y = 16'h1ff;
			16'h1b96: y = 16'h1ff;
			16'h1b97: y = 16'h1ff;
			16'h1b98: y = 16'h1ff;
			16'h1b99: y = 16'h1ff;
			16'h1b9a: y = 16'h1ff;
			16'h1b9b: y = 16'h1ff;
			16'h1b9c: y = 16'h1ff;
			16'h1b9d: y = 16'h1ff;
			16'h1b9e: y = 16'h1ff;
			16'h1b9f: y = 16'h1ff;
			16'h1ba0: y = 16'h1ff;
			16'h1ba1: y = 16'h1ff;
			16'h1ba2: y = 16'h1ff;
			16'h1ba3: y = 16'h1ff;
			16'h1ba4: y = 16'h1ff;
			16'h1ba5: y = 16'h1ff;
			16'h1ba6: y = 16'h1ff;
			16'h1ba7: y = 16'h1ff;
			16'h1ba8: y = 16'h1ff;
			16'h1ba9: y = 16'h1ff;
			16'h1baa: y = 16'h1ff;
			16'h1bab: y = 16'h1ff;
			16'h1bac: y = 16'h1ff;
			16'h1bad: y = 16'h1ff;
			16'h1bae: y = 16'h1ff;
			16'h1baf: y = 16'h1ff;
			16'h1bb0: y = 16'h1ff;
			16'h1bb1: y = 16'h1ff;
			16'h1bb2: y = 16'h1ff;
			16'h1bb3: y = 16'h1ff;
			16'h1bb4: y = 16'h1ff;
			16'h1bb5: y = 16'h1ff;
			16'h1bb6: y = 16'h1ff;
			16'h1bb7: y = 16'h1ff;
			16'h1bb8: y = 16'h1ff;
			16'h1bb9: y = 16'h1ff;
			16'h1bba: y = 16'h1ff;
			16'h1bbb: y = 16'h1ff;
			16'h1bbc: y = 16'h1ff;
			16'h1bbd: y = 16'h1ff;
			16'h1bbe: y = 16'h1ff;
			16'h1bbf: y = 16'h1ff;
			16'h1bc0: y = 16'h1ff;
			16'h1bc1: y = 16'h1ff;
			16'h1bc2: y = 16'h1ff;
			16'h1bc3: y = 16'h1ff;
			16'h1bc4: y = 16'h1ff;
			16'h1bc5: y = 16'h1ff;
			16'h1bc6: y = 16'h1ff;
			16'h1bc7: y = 16'h1ff;
			16'h1bc8: y = 16'h1ff;
			16'h1bc9: y = 16'h1ff;
			16'h1bca: y = 16'h1ff;
			16'h1bcb: y = 16'h1ff;
			16'h1bcc: y = 16'h1ff;
			16'h1bcd: y = 16'h1ff;
			16'h1bce: y = 16'h1ff;
			16'h1bcf: y = 16'h1ff;
			16'h1bd0: y = 16'h1ff;
			16'h1bd1: y = 16'h1ff;
			16'h1bd2: y = 16'h1ff;
			16'h1bd3: y = 16'h1ff;
			16'h1bd4: y = 16'h1ff;
			16'h1bd5: y = 16'h1ff;
			16'h1bd6: y = 16'h1ff;
			16'h1bd7: y = 16'h1ff;
			16'h1bd8: y = 16'h1ff;
			16'h1bd9: y = 16'h1ff;
			16'h1bda: y = 16'h1ff;
			16'h1bdb: y = 16'h1ff;
			16'h1bdc: y = 16'h1ff;
			16'h1bdd: y = 16'h1ff;
			16'h1bde: y = 16'h1ff;
			16'h1bdf: y = 16'h1ff;
			16'h1be0: y = 16'h1ff;
			16'h1be1: y = 16'h1ff;
			16'h1be2: y = 16'h1ff;
			16'h1be3: y = 16'h1ff;
			16'h1be4: y = 16'h1ff;
			16'h1be5: y = 16'h1ff;
			16'h1be6: y = 16'h1ff;
			16'h1be7: y = 16'h1ff;
			16'h1be8: y = 16'h1ff;
			16'h1be9: y = 16'h1ff;
			16'h1bea: y = 16'h1ff;
			16'h1beb: y = 16'h1ff;
			16'h1bec: y = 16'h1ff;
			16'h1bed: y = 16'h1ff;
			16'h1bee: y = 16'h1ff;
			16'h1bef: y = 16'h1ff;
			16'h1bf0: y = 16'h1ff;
			16'h1bf1: y = 16'h1ff;
			16'h1bf2: y = 16'h1ff;
			16'h1bf3: y = 16'h1ff;
			16'h1bf4: y = 16'h1ff;
			16'h1bf5: y = 16'h1ff;
			16'h1bf6: y = 16'h1ff;
			16'h1bf7: y = 16'h1ff;
			16'h1bf8: y = 16'h1ff;
			16'h1bf9: y = 16'h1ff;
			16'h1bfa: y = 16'h1ff;
			16'h1bfb: y = 16'h1ff;
			16'h1bfc: y = 16'h1ff;
			16'h1bfd: y = 16'h1ff;
			16'h1bfe: y = 16'h1ff;
			16'h1bff: y = 16'h1ff;
			16'h1c00: y = 16'h1ff;
			16'h1c01: y = 16'h1ff;
			16'h1c02: y = 16'h1ff;
			16'h1c03: y = 16'h1ff;
			16'h1c04: y = 16'h1ff;
			16'h1c05: y = 16'h1ff;
			16'h1c06: y = 16'h1ff;
			16'h1c07: y = 16'h1ff;
			16'h1c08: y = 16'h1ff;
			16'h1c09: y = 16'h1ff;
			16'h1c0a: y = 16'h1ff;
			16'h1c0b: y = 16'h1ff;
			16'h1c0c: y = 16'h1ff;
			16'h1c0d: y = 16'h1ff;
			16'h1c0e: y = 16'h1ff;
			16'h1c0f: y = 16'h1ff;
			16'h1c10: y = 16'h1ff;
			16'h1c11: y = 16'h1ff;
			16'h1c12: y = 16'h1ff;
			16'h1c13: y = 16'h1ff;
			16'h1c14: y = 16'h1ff;
			16'h1c15: y = 16'h1ff;
			16'h1c16: y = 16'h1ff;
			16'h1c17: y = 16'h1ff;
			16'h1c18: y = 16'h1ff;
			16'h1c19: y = 16'h1ff;
			16'h1c1a: y = 16'h1ff;
			16'h1c1b: y = 16'h1ff;
			16'h1c1c: y = 16'h1ff;
			16'h1c1d: y = 16'h1ff;
			16'h1c1e: y = 16'h1ff;
			16'h1c1f: y = 16'h1ff;
			16'h1c20: y = 16'h1ff;
			16'h1c21: y = 16'h1ff;
			16'h1c22: y = 16'h1ff;
			16'h1c23: y = 16'h1ff;
			16'h1c24: y = 16'h1ff;
			16'h1c25: y = 16'h1ff;
			16'h1c26: y = 16'h1ff;
			16'h1c27: y = 16'h1ff;
			16'h1c28: y = 16'h1ff;
			16'h1c29: y = 16'h1ff;
			16'h1c2a: y = 16'h1ff;
			16'h1c2b: y = 16'h1ff;
			16'h1c2c: y = 16'h1ff;
			16'h1c2d: y = 16'h1ff;
			16'h1c2e: y = 16'h1ff;
			16'h1c2f: y = 16'h1ff;
			16'h1c30: y = 16'h1ff;
			16'h1c31: y = 16'h1ff;
			16'h1c32: y = 16'h1ff;
			16'h1c33: y = 16'h1ff;
			16'h1c34: y = 16'h1ff;
			16'h1c35: y = 16'h1ff;
			16'h1c36: y = 16'h1ff;
			16'h1c37: y = 16'h1ff;
			16'h1c38: y = 16'h1ff;
			16'h1c39: y = 16'h1ff;
			16'h1c3a: y = 16'h1ff;
			16'h1c3b: y = 16'h1ff;
			16'h1c3c: y = 16'h1ff;
			16'h1c3d: y = 16'h1ff;
			16'h1c3e: y = 16'h1ff;
			16'h1c3f: y = 16'h1ff;
			16'h1c40: y = 16'h1ff;
			16'h1c41: y = 16'h1ff;
			16'h1c42: y = 16'h1ff;
			16'h1c43: y = 16'h1ff;
			16'h1c44: y = 16'h1ff;
			16'h1c45: y = 16'h1ff;
			16'h1c46: y = 16'h1ff;
			16'h1c47: y = 16'h1ff;
			16'h1c48: y = 16'h1ff;
			16'h1c49: y = 16'h1ff;
			16'h1c4a: y = 16'h1ff;
			16'h1c4b: y = 16'h1ff;
			16'h1c4c: y = 16'h1ff;
			16'h1c4d: y = 16'h1ff;
			16'h1c4e: y = 16'h1ff;
			16'h1c4f: y = 16'h1ff;
			16'h1c50: y = 16'h1ff;
			16'h1c51: y = 16'h1ff;
			16'h1c52: y = 16'h1ff;
			16'h1c53: y = 16'h1ff;
			16'h1c54: y = 16'h1ff;
			16'h1c55: y = 16'h1ff;
			16'h1c56: y = 16'h1ff;
			16'h1c57: y = 16'h1ff;
			16'h1c58: y = 16'h1ff;
			16'h1c59: y = 16'h1ff;
			16'h1c5a: y = 16'h1ff;
			16'h1c5b: y = 16'h1ff;
			16'h1c5c: y = 16'h1ff;
			16'h1c5d: y = 16'h1ff;
			16'h1c5e: y = 16'h1ff;
			16'h1c5f: y = 16'h1ff;
			16'h1c60: y = 16'h1ff;
			16'h1c61: y = 16'h1ff;
			16'h1c62: y = 16'h1ff;
			16'h1c63: y = 16'h1ff;
			16'h1c64: y = 16'h1ff;
			16'h1c65: y = 16'h1ff;
			16'h1c66: y = 16'h1ff;
			16'h1c67: y = 16'h1ff;
			16'h1c68: y = 16'h1ff;
			16'h1c69: y = 16'h1ff;
			16'h1c6a: y = 16'h1ff;
			16'h1c6b: y = 16'h1ff;
			16'h1c6c: y = 16'h1ff;
			16'h1c6d: y = 16'h1ff;
			16'h1c6e: y = 16'h1ff;
			16'h1c6f: y = 16'h1ff;
			16'h1c70: y = 16'h1ff;
			16'h1c71: y = 16'h1ff;
			16'h1c72: y = 16'h1ff;
			16'h1c73: y = 16'h1ff;
			16'h1c74: y = 16'h1ff;
			16'h1c75: y = 16'h1ff;
			16'h1c76: y = 16'h1ff;
			16'h1c77: y = 16'h1ff;
			16'h1c78: y = 16'h1ff;
			16'h1c79: y = 16'h1ff;
			16'h1c7a: y = 16'h1ff;
			16'h1c7b: y = 16'h1ff;
			16'h1c7c: y = 16'h1ff;
			16'h1c7d: y = 16'h1ff;
			16'h1c7e: y = 16'h1ff;
			16'h1c7f: y = 16'h1ff;
			16'h1c80: y = 16'h1ff;
			16'h1c81: y = 16'h1ff;
			16'h1c82: y = 16'h1ff;
			16'h1c83: y = 16'h1ff;
			16'h1c84: y = 16'h1ff;
			16'h1c85: y = 16'h1ff;
			16'h1c86: y = 16'h1ff;
			16'h1c87: y = 16'h1ff;
			16'h1c88: y = 16'h1ff;
			16'h1c89: y = 16'h1ff;
			16'h1c8a: y = 16'h1ff;
			16'h1c8b: y = 16'h1ff;
			16'h1c8c: y = 16'h1ff;
			16'h1c8d: y = 16'h1ff;
			16'h1c8e: y = 16'h1ff;
			16'h1c8f: y = 16'h1ff;
			16'h1c90: y = 16'h1ff;
			16'h1c91: y = 16'h1ff;
			16'h1c92: y = 16'h1ff;
			16'h1c93: y = 16'h1ff;
			16'h1c94: y = 16'h1ff;
			16'h1c95: y = 16'h1ff;
			16'h1c96: y = 16'h1ff;
			16'h1c97: y = 16'h1ff;
			16'h1c98: y = 16'h1ff;
			16'h1c99: y = 16'h1ff;
			16'h1c9a: y = 16'h1ff;
			16'h1c9b: y = 16'h1ff;
			16'h1c9c: y = 16'h1ff;
			16'h1c9d: y = 16'h1ff;
			16'h1c9e: y = 16'h1ff;
			16'h1c9f: y = 16'h1ff;
			16'h1ca0: y = 16'h1ff;
			16'h1ca1: y = 16'h1ff;
			16'h1ca2: y = 16'h1ff;
			16'h1ca3: y = 16'h1ff;
			16'h1ca4: y = 16'h1ff;
			16'h1ca5: y = 16'h1ff;
			16'h1ca6: y = 16'h1ff;
			16'h1ca7: y = 16'h1ff;
			16'h1ca8: y = 16'h1ff;
			16'h1ca9: y = 16'h1ff;
			16'h1caa: y = 16'h1ff;
			16'h1cab: y = 16'h1ff;
			16'h1cac: y = 16'h1ff;
			16'h1cad: y = 16'h1ff;
			16'h1cae: y = 16'h1ff;
			16'h1caf: y = 16'h1ff;
			16'h1cb0: y = 16'h1ff;
			16'h1cb1: y = 16'h1ff;
			16'h1cb2: y = 16'h1ff;
			16'h1cb3: y = 16'h1ff;
			16'h1cb4: y = 16'h1ff;
			16'h1cb5: y = 16'h1ff;
			16'h1cb6: y = 16'h1ff;
			16'h1cb7: y = 16'h1ff;
			16'h1cb8: y = 16'h1ff;
			16'h1cb9: y = 16'h1ff;
			16'h1cba: y = 16'h1ff;
			16'h1cbb: y = 16'h1ff;
			16'h1cbc: y = 16'h1ff;
			16'h1cbd: y = 16'h1ff;
			16'h1cbe: y = 16'h1ff;
			16'h1cbf: y = 16'h1ff;
			16'h1cc0: y = 16'h1ff;
			16'h1cc1: y = 16'h1ff;
			16'h1cc2: y = 16'h1ff;
			16'h1cc3: y = 16'h1ff;
			16'h1cc4: y = 16'h1ff;
			16'h1cc5: y = 16'h1ff;
			16'h1cc6: y = 16'h1ff;
			16'h1cc7: y = 16'h1ff;
			16'h1cc8: y = 16'h1ff;
			16'h1cc9: y = 16'h1ff;
			16'h1cca: y = 16'h1ff;
			16'h1ccb: y = 16'h1ff;
			16'h1ccc: y = 16'h1ff;
			16'h1ccd: y = 16'h1ff;
			16'h1cce: y = 16'h1ff;
			16'h1ccf: y = 16'h1ff;
			16'h1cd0: y = 16'h1ff;
			16'h1cd1: y = 16'h1ff;
			16'h1cd2: y = 16'h1ff;
			16'h1cd3: y = 16'h1ff;
			16'h1cd4: y = 16'h1ff;
			16'h1cd5: y = 16'h1ff;
			16'h1cd6: y = 16'h1ff;
			16'h1cd7: y = 16'h1ff;
			16'h1cd8: y = 16'h1ff;
			16'h1cd9: y = 16'h1ff;
			16'h1cda: y = 16'h1ff;
			16'h1cdb: y = 16'h1ff;
			16'h1cdc: y = 16'h1ff;
			16'h1cdd: y = 16'h1ff;
			16'h1cde: y = 16'h1ff;
			16'h1cdf: y = 16'h1ff;
			16'h1ce0: y = 16'h1ff;
			16'h1ce1: y = 16'h1ff;
			16'h1ce2: y = 16'h1ff;
			16'h1ce3: y = 16'h1ff;
			16'h1ce4: y = 16'h1ff;
			16'h1ce5: y = 16'h1ff;
			16'h1ce6: y = 16'h1ff;
			16'h1ce7: y = 16'h1ff;
			16'h1ce8: y = 16'h1ff;
			16'h1ce9: y = 16'h1ff;
			16'h1cea: y = 16'h1ff;
			16'h1ceb: y = 16'h1ff;
			16'h1cec: y = 16'h1ff;
			16'h1ced: y = 16'h1ff;
			16'h1cee: y = 16'h1ff;
			16'h1cef: y = 16'h1ff;
			16'h1cf0: y = 16'h1ff;
			16'h1cf1: y = 16'h1ff;
			16'h1cf2: y = 16'h1ff;
			16'h1cf3: y = 16'h1ff;
			16'h1cf4: y = 16'h1ff;
			16'h1cf5: y = 16'h1ff;
			16'h1cf6: y = 16'h1ff;
			16'h1cf7: y = 16'h1ff;
			16'h1cf8: y = 16'h1ff;
			16'h1cf9: y = 16'h1ff;
			16'h1cfa: y = 16'h1ff;
			16'h1cfb: y = 16'h1ff;
			16'h1cfc: y = 16'h1ff;
			16'h1cfd: y = 16'h1ff;
			16'h1cfe: y = 16'h1ff;
			16'h1cff: y = 16'h1ff;
			16'h1d00: y = 16'h1ff;
			16'h1d01: y = 16'h1ff;
			16'h1d02: y = 16'h1ff;
			16'h1d03: y = 16'h1ff;
			16'h1d04: y = 16'h1ff;
			16'h1d05: y = 16'h1ff;
			16'h1d06: y = 16'h1ff;
			16'h1d07: y = 16'h1ff;
			16'h1d08: y = 16'h1ff;
			16'h1d09: y = 16'h1ff;
			16'h1d0a: y = 16'h1ff;
			16'h1d0b: y = 16'h1ff;
			16'h1d0c: y = 16'h1ff;
			16'h1d0d: y = 16'h1ff;
			16'h1d0e: y = 16'h1ff;
			16'h1d0f: y = 16'h1ff;
			16'h1d10: y = 16'h1ff;
			16'h1d11: y = 16'h1ff;
			16'h1d12: y = 16'h1ff;
			16'h1d13: y = 16'h1ff;
			16'h1d14: y = 16'h1ff;
			16'h1d15: y = 16'h1ff;
			16'h1d16: y = 16'h1ff;
			16'h1d17: y = 16'h1ff;
			16'h1d18: y = 16'h1ff;
			16'h1d19: y = 16'h1ff;
			16'h1d1a: y = 16'h1ff;
			16'h1d1b: y = 16'h1ff;
			16'h1d1c: y = 16'h1ff;
			16'h1d1d: y = 16'h1ff;
			16'h1d1e: y = 16'h1ff;
			16'h1d1f: y = 16'h1ff;
			16'h1d20: y = 16'h1ff;
			16'h1d21: y = 16'h1ff;
			16'h1d22: y = 16'h1ff;
			16'h1d23: y = 16'h1ff;
			16'h1d24: y = 16'h1ff;
			16'h1d25: y = 16'h1ff;
			16'h1d26: y = 16'h1ff;
			16'h1d27: y = 16'h1ff;
			16'h1d28: y = 16'h1ff;
			16'h1d29: y = 16'h1ff;
			16'h1d2a: y = 16'h1ff;
			16'h1d2b: y = 16'h1ff;
			16'h1d2c: y = 16'h1ff;
			16'h1d2d: y = 16'h1ff;
			16'h1d2e: y = 16'h1ff;
			16'h1d2f: y = 16'h1ff;
			16'h1d30: y = 16'h1ff;
			16'h1d31: y = 16'h1ff;
			16'h1d32: y = 16'h1ff;
			16'h1d33: y = 16'h1ff;
			16'h1d34: y = 16'h1ff;
			16'h1d35: y = 16'h1ff;
			16'h1d36: y = 16'h1ff;
			16'h1d37: y = 16'h1ff;
			16'h1d38: y = 16'h1ff;
			16'h1d39: y = 16'h1ff;
			16'h1d3a: y = 16'h1ff;
			16'h1d3b: y = 16'h1ff;
			16'h1d3c: y = 16'h1ff;
			16'h1d3d: y = 16'h1ff;
			16'h1d3e: y = 16'h1ff;
			16'h1d3f: y = 16'h1ff;
			16'h1d40: y = 16'h1ff;
			16'h1d41: y = 16'h1ff;
			16'h1d42: y = 16'h1ff;
			16'h1d43: y = 16'h1ff;
			16'h1d44: y = 16'h1ff;
			16'h1d45: y = 16'h1ff;
			16'h1d46: y = 16'h1ff;
			16'h1d47: y = 16'h1ff;
			16'h1d48: y = 16'h1ff;
			16'h1d49: y = 16'h1ff;
			16'h1d4a: y = 16'h1ff;
			16'h1d4b: y = 16'h1ff;
			16'h1d4c: y = 16'h1ff;
			16'h1d4d: y = 16'h1ff;
			16'h1d4e: y = 16'h1ff;
			16'h1d4f: y = 16'h1ff;
			16'h1d50: y = 16'h1ff;
			16'h1d51: y = 16'h1ff;
			16'h1d52: y = 16'h1ff;
			16'h1d53: y = 16'h1ff;
			16'h1d54: y = 16'h1ff;
			16'h1d55: y = 16'h1ff;
			16'h1d56: y = 16'h1ff;
			16'h1d57: y = 16'h1ff;
			16'h1d58: y = 16'h1ff;
			16'h1d59: y = 16'h1ff;
			16'h1d5a: y = 16'h1ff;
			16'h1d5b: y = 16'h1ff;
			16'h1d5c: y = 16'h1ff;
			16'h1d5d: y = 16'h1ff;
			16'h1d5e: y = 16'h1ff;
			16'h1d5f: y = 16'h1ff;
			16'h1d60: y = 16'h1ff;
			16'h1d61: y = 16'h1ff;
			16'h1d62: y = 16'h1ff;
			16'h1d63: y = 16'h1ff;
			16'h1d64: y = 16'h1ff;
			16'h1d65: y = 16'h1ff;
			16'h1d66: y = 16'h1ff;
			16'h1d67: y = 16'h1ff;
			16'h1d68: y = 16'h1ff;
			16'h1d69: y = 16'h1ff;
			16'h1d6a: y = 16'h1ff;
			16'h1d6b: y = 16'h1ff;
			16'h1d6c: y = 16'h1ff;
			16'h1d6d: y = 16'h1ff;
			16'h1d6e: y = 16'h1ff;
			16'h1d6f: y = 16'h1ff;
			16'h1d70: y = 16'h1ff;
			16'h1d71: y = 16'h1ff;
			16'h1d72: y = 16'h1ff;
			16'h1d73: y = 16'h1ff;
			16'h1d74: y = 16'h1ff;
			16'h1d75: y = 16'h1ff;
			16'h1d76: y = 16'h1ff;
			16'h1d77: y = 16'h1ff;
			16'h1d78: y = 16'h1ff;
			16'h1d79: y = 16'h1ff;
			16'h1d7a: y = 16'h1ff;
			16'h1d7b: y = 16'h1ff;
			16'h1d7c: y = 16'h1ff;
			16'h1d7d: y = 16'h1ff;
			16'h1d7e: y = 16'h1ff;
			16'h1d7f: y = 16'h1ff;
			16'h1d80: y = 16'h1ff;
			16'h1d81: y = 16'h1ff;
			16'h1d82: y = 16'h1ff;
			16'h1d83: y = 16'h1ff;
			16'h1d84: y = 16'h1ff;
			16'h1d85: y = 16'h1ff;
			16'h1d86: y = 16'h1ff;
			16'h1d87: y = 16'h1ff;
			16'h1d88: y = 16'h1ff;
			16'h1d89: y = 16'h1ff;
			16'h1d8a: y = 16'h1ff;
			16'h1d8b: y = 16'h1ff;
			16'h1d8c: y = 16'h1ff;
			16'h1d8d: y = 16'h1ff;
			16'h1d8e: y = 16'h1ff;
			16'h1d8f: y = 16'h1ff;
			16'h1d90: y = 16'h1ff;
			16'h1d91: y = 16'h1ff;
			16'h1d92: y = 16'h1ff;
			16'h1d93: y = 16'h1ff;
			16'h1d94: y = 16'h1ff;
			16'h1d95: y = 16'h1ff;
			16'h1d96: y = 16'h1ff;
			16'h1d97: y = 16'h1ff;
			16'h1d98: y = 16'h1ff;
			16'h1d99: y = 16'h1ff;
			16'h1d9a: y = 16'h1ff;
			16'h1d9b: y = 16'h1ff;
			16'h1d9c: y = 16'h1ff;
			16'h1d9d: y = 16'h1ff;
			16'h1d9e: y = 16'h1ff;
			16'h1d9f: y = 16'h1ff;
			16'h1da0: y = 16'h1ff;
			16'h1da1: y = 16'h1ff;
			16'h1da2: y = 16'h1ff;
			16'h1da3: y = 16'h1ff;
			16'h1da4: y = 16'h1ff;
			16'h1da5: y = 16'h1ff;
			16'h1da6: y = 16'h1ff;
			16'h1da7: y = 16'h1ff;
			16'h1da8: y = 16'h1ff;
			16'h1da9: y = 16'h1ff;
			16'h1daa: y = 16'h1ff;
			16'h1dab: y = 16'h1ff;
			16'h1dac: y = 16'h1ff;
			16'h1dad: y = 16'h1ff;
			16'h1dae: y = 16'h1ff;
			16'h1daf: y = 16'h1ff;
			16'h1db0: y = 16'h1ff;
			16'h1db1: y = 16'h1ff;
			16'h1db2: y = 16'h1ff;
			16'h1db3: y = 16'h1ff;
			16'h1db4: y = 16'h1ff;
			16'h1db5: y = 16'h1ff;
			16'h1db6: y = 16'h1ff;
			16'h1db7: y = 16'h1ff;
			16'h1db8: y = 16'h1ff;
			16'h1db9: y = 16'h1ff;
			16'h1dba: y = 16'h1ff;
			16'h1dbb: y = 16'h1ff;
			16'h1dbc: y = 16'h1ff;
			16'h1dbd: y = 16'h1ff;
			16'h1dbe: y = 16'h1ff;
			16'h1dbf: y = 16'h1ff;
			16'h1dc0: y = 16'h1ff;
			16'h1dc1: y = 16'h1ff;
			16'h1dc2: y = 16'h1ff;
			16'h1dc3: y = 16'h1ff;
			16'h1dc4: y = 16'h1ff;
			16'h1dc5: y = 16'h1ff;
			16'h1dc6: y = 16'h1ff;
			16'h1dc7: y = 16'h1ff;
			16'h1dc8: y = 16'h1ff;
			16'h1dc9: y = 16'h1ff;
			16'h1dca: y = 16'h1ff;
			16'h1dcb: y = 16'h1ff;
			16'h1dcc: y = 16'h1ff;
			16'h1dcd: y = 16'h1ff;
			16'h1dce: y = 16'h1ff;
			16'h1dcf: y = 16'h1ff;
			16'h1dd0: y = 16'h1ff;
			16'h1dd1: y = 16'h1ff;
			16'h1dd2: y = 16'h1ff;
			16'h1dd3: y = 16'h1ff;
			16'h1dd4: y = 16'h1ff;
			16'h1dd5: y = 16'h1ff;
			16'h1dd6: y = 16'h1ff;
			16'h1dd7: y = 16'h1ff;
			16'h1dd8: y = 16'h1ff;
			16'h1dd9: y = 16'h1ff;
			16'h1dda: y = 16'h1ff;
			16'h1ddb: y = 16'h1ff;
			16'h1ddc: y = 16'h1ff;
			16'h1ddd: y = 16'h1ff;
			16'h1dde: y = 16'h1ff;
			16'h1ddf: y = 16'h1ff;
			16'h1de0: y = 16'h1ff;
			16'h1de1: y = 16'h1ff;
			16'h1de2: y = 16'h1ff;
			16'h1de3: y = 16'h1ff;
			16'h1de4: y = 16'h1ff;
			16'h1de5: y = 16'h1ff;
			16'h1de6: y = 16'h1ff;
			16'h1de7: y = 16'h1ff;
			16'h1de8: y = 16'h1ff;
			16'h1de9: y = 16'h1ff;
			16'h1dea: y = 16'h1ff;
			16'h1deb: y = 16'h1ff;
			16'h1dec: y = 16'h1ff;
			16'h1ded: y = 16'h1ff;
			16'h1dee: y = 16'h1ff;
			16'h1def: y = 16'h1ff;
			16'h1df0: y = 16'h1ff;
			16'h1df1: y = 16'h1ff;
			16'h1df2: y = 16'h1ff;
			16'h1df3: y = 16'h1ff;
			16'h1df4: y = 16'h1ff;
			16'h1df5: y = 16'h1ff;
			16'h1df6: y = 16'h1ff;
			16'h1df7: y = 16'h1ff;
			16'h1df8: y = 16'h1ff;
			16'h1df9: y = 16'h1ff;
			16'h1dfa: y = 16'h1ff;
			16'h1dfb: y = 16'h1ff;
			16'h1dfc: y = 16'h1ff;
			16'h1dfd: y = 16'h1ff;
			16'h1dfe: y = 16'h1ff;
			16'h1dff: y = 16'h1ff;
			16'h1e00: y = 16'h1ff;
			16'h1e01: y = 16'h1ff;
			16'h1e02: y = 16'h1ff;
			16'h1e03: y = 16'h1ff;
			16'h1e04: y = 16'h1ff;
			16'h1e05: y = 16'h1ff;
			16'h1e06: y = 16'h1ff;
			16'h1e07: y = 16'h1ff;
			16'h1e08: y = 16'h1ff;
			16'h1e09: y = 16'h1ff;
			16'h1e0a: y = 16'h1ff;
			16'h1e0b: y = 16'h1ff;
			16'h1e0c: y = 16'h1ff;
			16'h1e0d: y = 16'h1ff;
			16'h1e0e: y = 16'h1ff;
			16'h1e0f: y = 16'h1ff;
			16'h1e10: y = 16'h1ff;
			16'h1e11: y = 16'h1ff;
			16'h1e12: y = 16'h1ff;
			16'h1e13: y = 16'h1ff;
			16'h1e14: y = 16'h1ff;
			16'h1e15: y = 16'h1ff;
			16'h1e16: y = 16'h1ff;
			16'h1e17: y = 16'h1ff;
			16'h1e18: y = 16'h1ff;
			16'h1e19: y = 16'h1ff;
			16'h1e1a: y = 16'h1ff;
			16'h1e1b: y = 16'h1ff;
			16'h1e1c: y = 16'h1ff;
			16'h1e1d: y = 16'h1ff;
			16'h1e1e: y = 16'h1ff;
			16'h1e1f: y = 16'h1ff;
			16'h1e20: y = 16'h1ff;
			16'h1e21: y = 16'h1ff;
			16'h1e22: y = 16'h1ff;
			16'h1e23: y = 16'h1ff;
			16'h1e24: y = 16'h1ff;
			16'h1e25: y = 16'h1ff;
			16'h1e26: y = 16'h1ff;
			16'h1e27: y = 16'h1ff;
			16'h1e28: y = 16'h1ff;
			16'h1e29: y = 16'h1ff;
			16'h1e2a: y = 16'h1ff;
			16'h1e2b: y = 16'h1ff;
			16'h1e2c: y = 16'h1ff;
			16'h1e2d: y = 16'h1ff;
			16'h1e2e: y = 16'h1ff;
			16'h1e2f: y = 16'h1ff;
			16'h1e30: y = 16'h1ff;
			16'h1e31: y = 16'h1ff;
			16'h1e32: y = 16'h1ff;
			16'h1e33: y = 16'h1ff;
			16'h1e34: y = 16'h1ff;
			16'h1e35: y = 16'h1ff;
			16'h1e36: y = 16'h1ff;
			16'h1e37: y = 16'h1ff;
			16'h1e38: y = 16'h1ff;
			16'h1e39: y = 16'h1ff;
			16'h1e3a: y = 16'h1ff;
			16'h1e3b: y = 16'h1ff;
			16'h1e3c: y = 16'h1ff;
			16'h1e3d: y = 16'h1ff;
			16'h1e3e: y = 16'h1ff;
			16'h1e3f: y = 16'h1ff;
			16'h1e40: y = 16'h1ff;
			16'h1e41: y = 16'h1ff;
			16'h1e42: y = 16'h1ff;
			16'h1e43: y = 16'h1ff;
			16'h1e44: y = 16'h1ff;
			16'h1e45: y = 16'h1ff;
			16'h1e46: y = 16'h1ff;
			16'h1e47: y = 16'h1ff;
			16'h1e48: y = 16'h1ff;
			16'h1e49: y = 16'h1ff;
			16'h1e4a: y = 16'h1ff;
			16'h1e4b: y = 16'h1ff;
			16'h1e4c: y = 16'h1ff;
			16'h1e4d: y = 16'h1ff;
			16'h1e4e: y = 16'h1ff;
			16'h1e4f: y = 16'h1ff;
			16'h1e50: y = 16'h1ff;
			16'h1e51: y = 16'h1ff;
			16'h1e52: y = 16'h1ff;
			16'h1e53: y = 16'h1ff;
			16'h1e54: y = 16'h1ff;
			16'h1e55: y = 16'h1ff;
			16'h1e56: y = 16'h1ff;
			16'h1e57: y = 16'h1ff;
			16'h1e58: y = 16'h1ff;
			16'h1e59: y = 16'h1ff;
			16'h1e5a: y = 16'h1ff;
			16'h1e5b: y = 16'h1ff;
			16'h1e5c: y = 16'h1ff;
			16'h1e5d: y = 16'h1ff;
			16'h1e5e: y = 16'h1ff;
			16'h1e5f: y = 16'h1ff;
			16'h1e60: y = 16'h1ff;
			16'h1e61: y = 16'h1ff;
			16'h1e62: y = 16'h1ff;
			16'h1e63: y = 16'h1ff;
			16'h1e64: y = 16'h1ff;
			16'h1e65: y = 16'h1ff;
			16'h1e66: y = 16'h1ff;
			16'h1e67: y = 16'h1ff;
			16'h1e68: y = 16'h1ff;
			16'h1e69: y = 16'h1ff;
			16'h1e6a: y = 16'h1ff;
			16'h1e6b: y = 16'h1ff;
			16'h1e6c: y = 16'h1ff;
			16'h1e6d: y = 16'h1ff;
			16'h1e6e: y = 16'h1ff;
			16'h1e6f: y = 16'h1ff;
			16'h1e70: y = 16'h1ff;
			16'h1e71: y = 16'h1ff;
			16'h1e72: y = 16'h1ff;
			16'h1e73: y = 16'h1ff;
			16'h1e74: y = 16'h1ff;
			16'h1e75: y = 16'h1ff;
			16'h1e76: y = 16'h1ff;
			16'h1e77: y = 16'h1ff;
			16'h1e78: y = 16'h1ff;
			16'h1e79: y = 16'h1ff;
			16'h1e7a: y = 16'h1ff;
			16'h1e7b: y = 16'h1ff;
			16'h1e7c: y = 16'h1ff;
			16'h1e7d: y = 16'h1ff;
			16'h1e7e: y = 16'h1ff;
			16'h1e7f: y = 16'h1ff;
			16'h1e80: y = 16'h1ff;
			16'h1e81: y = 16'h1ff;
			16'h1e82: y = 16'h1ff;
			16'h1e83: y = 16'h1ff;
			16'h1e84: y = 16'h1ff;
			16'h1e85: y = 16'h1ff;
			16'h1e86: y = 16'h1ff;
			16'h1e87: y = 16'h1ff;
			16'h1e88: y = 16'h1ff;
			16'h1e89: y = 16'h1ff;
			16'h1e8a: y = 16'h1ff;
			16'h1e8b: y = 16'h1ff;
			16'h1e8c: y = 16'h1ff;
			16'h1e8d: y = 16'h1ff;
			16'h1e8e: y = 16'h1ff;
			16'h1e8f: y = 16'h1ff;
			16'h1e90: y = 16'h1ff;
			16'h1e91: y = 16'h1ff;
			16'h1e92: y = 16'h1ff;
			16'h1e93: y = 16'h1ff;
			16'h1e94: y = 16'h1ff;
			16'h1e95: y = 16'h1ff;
			16'h1e96: y = 16'h1ff;
			16'h1e97: y = 16'h1ff;
			16'h1e98: y = 16'h1ff;
			16'h1e99: y = 16'h1ff;
			16'h1e9a: y = 16'h1ff;
			16'h1e9b: y = 16'h1ff;
			16'h1e9c: y = 16'h1ff;
			16'h1e9d: y = 16'h1ff;
			16'h1e9e: y = 16'h1ff;
			16'h1e9f: y = 16'h1ff;
			16'h1ea0: y = 16'h1ff;
			16'h1ea1: y = 16'h1ff;
			16'h1ea2: y = 16'h1ff;
			16'h1ea3: y = 16'h1ff;
			16'h1ea4: y = 16'h1ff;
			16'h1ea5: y = 16'h1ff;
			16'h1ea6: y = 16'h1ff;
			16'h1ea7: y = 16'h1ff;
			16'h1ea8: y = 16'h1ff;
			16'h1ea9: y = 16'h1ff;
			16'h1eaa: y = 16'h1ff;
			16'h1eab: y = 16'h1ff;
			16'h1eac: y = 16'h1ff;
			16'h1ead: y = 16'h1ff;
			16'h1eae: y = 16'h1ff;
			16'h1eaf: y = 16'h1ff;
			16'h1eb0: y = 16'h1ff;
			16'h1eb1: y = 16'h1ff;
			16'h1eb2: y = 16'h1ff;
			16'h1eb3: y = 16'h1ff;
			16'h1eb4: y = 16'h1ff;
			16'h1eb5: y = 16'h1ff;
			16'h1eb6: y = 16'h1ff;
			16'h1eb7: y = 16'h1ff;
			16'h1eb8: y = 16'h1ff;
			16'h1eb9: y = 16'h1ff;
			16'h1eba: y = 16'h1ff;
			16'h1ebb: y = 16'h1ff;
			16'h1ebc: y = 16'h1ff;
			16'h1ebd: y = 16'h1ff;
			16'h1ebe: y = 16'h1ff;
			16'h1ebf: y = 16'h1ff;
			16'h1ec0: y = 16'h1ff;
			16'h1ec1: y = 16'h1ff;
			16'h1ec2: y = 16'h1ff;
			16'h1ec3: y = 16'h1ff;
			16'h1ec4: y = 16'h1ff;
			16'h1ec5: y = 16'h1ff;
			16'h1ec6: y = 16'h1ff;
			16'h1ec7: y = 16'h1ff;
			16'h1ec8: y = 16'h1ff;
			16'h1ec9: y = 16'h1ff;
			16'h1eca: y = 16'h1ff;
			16'h1ecb: y = 16'h1ff;
			16'h1ecc: y = 16'h1ff;
			16'h1ecd: y = 16'h1ff;
			16'h1ece: y = 16'h1ff;
			16'h1ecf: y = 16'h1ff;
			16'h1ed0: y = 16'h1ff;
			16'h1ed1: y = 16'h1ff;
			16'h1ed2: y = 16'h1ff;
			16'h1ed3: y = 16'h1ff;
			16'h1ed4: y = 16'h1ff;
			16'h1ed5: y = 16'h1ff;
			16'h1ed6: y = 16'h1ff;
			16'h1ed7: y = 16'h1ff;
			16'h1ed8: y = 16'h1ff;
			16'h1ed9: y = 16'h1ff;
			16'h1eda: y = 16'h1ff;
			16'h1edb: y = 16'h1ff;
			16'h1edc: y = 16'h1ff;
			16'h1edd: y = 16'h1ff;
			16'h1ede: y = 16'h1ff;
			16'h1edf: y = 16'h1ff;
			16'h1ee0: y = 16'h1ff;
			16'h1ee1: y = 16'h1ff;
			16'h1ee2: y = 16'h1ff;
			16'h1ee3: y = 16'h1ff;
			16'h1ee4: y = 16'h1ff;
			16'h1ee5: y = 16'h1ff;
			16'h1ee6: y = 16'h1ff;
			16'h1ee7: y = 16'h1ff;
			16'h1ee8: y = 16'h1ff;
			16'h1ee9: y = 16'h1ff;
			16'h1eea: y = 16'h1ff;
			16'h1eeb: y = 16'h1ff;
			16'h1eec: y = 16'h1ff;
			16'h1eed: y = 16'h1ff;
			16'h1eee: y = 16'h1ff;
			16'h1eef: y = 16'h1ff;
			16'h1ef0: y = 16'h1ff;
			16'h1ef1: y = 16'h1ff;
			16'h1ef2: y = 16'h1ff;
			16'h1ef3: y = 16'h1ff;
			16'h1ef4: y = 16'h1ff;
			16'h1ef5: y = 16'h1ff;
			16'h1ef6: y = 16'h1ff;
			16'h1ef7: y = 16'h1ff;
			16'h1ef8: y = 16'h1ff;
			16'h1ef9: y = 16'h1ff;
			16'h1efa: y = 16'h1ff;
			16'h1efb: y = 16'h1ff;
			16'h1efc: y = 16'h1ff;
			16'h1efd: y = 16'h1ff;
			16'h1efe: y = 16'h1ff;
			16'h1eff: y = 16'h1ff;
			16'h1f00: y = 16'h1ff;
			16'h1f01: y = 16'h1ff;
			16'h1f02: y = 16'h1ff;
			16'h1f03: y = 16'h1ff;
			16'h1f04: y = 16'h1ff;
			16'h1f05: y = 16'h1ff;
			16'h1f06: y = 16'h1ff;
			16'h1f07: y = 16'h1ff;
			16'h1f08: y = 16'h1ff;
			16'h1f09: y = 16'h1ff;
			16'h1f0a: y = 16'h1ff;
			16'h1f0b: y = 16'h1ff;
			16'h1f0c: y = 16'h1ff;
			16'h1f0d: y = 16'h1ff;
			16'h1f0e: y = 16'h1ff;
			16'h1f0f: y = 16'h1ff;
			16'h1f10: y = 16'h1ff;
			16'h1f11: y = 16'h1ff;
			16'h1f12: y = 16'h1ff;
			16'h1f13: y = 16'h1ff;
			16'h1f14: y = 16'h1ff;
			16'h1f15: y = 16'h1ff;
			16'h1f16: y = 16'h1ff;
			16'h1f17: y = 16'h1ff;
			16'h1f18: y = 16'h1ff;
			16'h1f19: y = 16'h1ff;
			16'h1f1a: y = 16'h1ff;
			16'h1f1b: y = 16'h1ff;
			16'h1f1c: y = 16'h1ff;
			16'h1f1d: y = 16'h1ff;
			16'h1f1e: y = 16'h1ff;
			16'h1f1f: y = 16'h1ff;
			16'h1f20: y = 16'h1ff;
			16'h1f21: y = 16'h1ff;
			16'h1f22: y = 16'h1ff;
			16'h1f23: y = 16'h1ff;
			16'h1f24: y = 16'h1ff;
			16'h1f25: y = 16'h1ff;
			16'h1f26: y = 16'h1ff;
			16'h1f27: y = 16'h1ff;
			16'h1f28: y = 16'h1ff;
			16'h1f29: y = 16'h1ff;
			16'h1f2a: y = 16'h1ff;
			16'h1f2b: y = 16'h1ff;
			16'h1f2c: y = 16'h1ff;
			16'h1f2d: y = 16'h1ff;
			16'h1f2e: y = 16'h1ff;
			16'h1f2f: y = 16'h1ff;
			16'h1f30: y = 16'h1ff;
			16'h1f31: y = 16'h1ff;
			16'h1f32: y = 16'h1ff;
			16'h1f33: y = 16'h1ff;
			16'h1f34: y = 16'h1ff;
			16'h1f35: y = 16'h1ff;
			16'h1f36: y = 16'h1ff;
			16'h1f37: y = 16'h1ff;
			16'h1f38: y = 16'h1ff;
			16'h1f39: y = 16'h1ff;
			16'h1f3a: y = 16'h1ff;
			16'h1f3b: y = 16'h1ff;
			16'h1f3c: y = 16'h1ff;
			16'h1f3d: y = 16'h1ff;
			16'h1f3e: y = 16'h1ff;
			16'h1f3f: y = 16'h1ff;
			16'h1f40: y = 16'h1ff;
			16'h1f41: y = 16'h1ff;
			16'h1f42: y = 16'h1ff;
			16'h1f43: y = 16'h1ff;
			16'h1f44: y = 16'h1ff;
			16'h1f45: y = 16'h1ff;
			16'h1f46: y = 16'h1ff;
			16'h1f47: y = 16'h1ff;
			16'h1f48: y = 16'h1ff;
			16'h1f49: y = 16'h1ff;
			16'h1f4a: y = 16'h1ff;
			16'h1f4b: y = 16'h1ff;
			16'h1f4c: y = 16'h1ff;
			16'h1f4d: y = 16'h1ff;
			16'h1f4e: y = 16'h1ff;
			16'h1f4f: y = 16'h1ff;
			16'h1f50: y = 16'h1ff;
			16'h1f51: y = 16'h1ff;
			16'h1f52: y = 16'h1ff;
			16'h1f53: y = 16'h1ff;
			16'h1f54: y = 16'h1ff;
			16'h1f55: y = 16'h1ff;
			16'h1f56: y = 16'h1ff;
			16'h1f57: y = 16'h1ff;
			16'h1f58: y = 16'h1ff;
			16'h1f59: y = 16'h1ff;
			16'h1f5a: y = 16'h1ff;
			16'h1f5b: y = 16'h1ff;
			16'h1f5c: y = 16'h1ff;
			16'h1f5d: y = 16'h1ff;
			16'h1f5e: y = 16'h1ff;
			16'h1f5f: y = 16'h1ff;
			16'h1f60: y = 16'h1ff;
			16'h1f61: y = 16'h1ff;
			16'h1f62: y = 16'h1ff;
			16'h1f63: y = 16'h1ff;
			16'h1f64: y = 16'h1ff;
			16'h1f65: y = 16'h1ff;
			16'h1f66: y = 16'h1ff;
			16'h1f67: y = 16'h1ff;
			16'h1f68: y = 16'h1ff;
			16'h1f69: y = 16'h1ff;
			16'h1f6a: y = 16'h1ff;
			16'h1f6b: y = 16'h1ff;
			16'h1f6c: y = 16'h1ff;
			16'h1f6d: y = 16'h1ff;
			16'h1f6e: y = 16'h1ff;
			16'h1f6f: y = 16'h1ff;
			16'h1f70: y = 16'h1ff;
			16'h1f71: y = 16'h1ff;
			16'h1f72: y = 16'h1ff;
			16'h1f73: y = 16'h1ff;
			16'h1f74: y = 16'h1ff;
			16'h1f75: y = 16'h1ff;
			16'h1f76: y = 16'h1ff;
			16'h1f77: y = 16'h1ff;
			16'h1f78: y = 16'h1ff;
			16'h1f79: y = 16'h1ff;
			16'h1f7a: y = 16'h1ff;
			16'h1f7b: y = 16'h1ff;
			16'h1f7c: y = 16'h1ff;
			16'h1f7d: y = 16'h1ff;
			16'h1f7e: y = 16'h1ff;
			16'h1f7f: y = 16'h1ff;
			16'h1f80: y = 16'h1ff;
			16'h1f81: y = 16'h1ff;
			16'h1f82: y = 16'h1ff;
			16'h1f83: y = 16'h1ff;
			16'h1f84: y = 16'h1ff;
			16'h1f85: y = 16'h1ff;
			16'h1f86: y = 16'h1ff;
			16'h1f87: y = 16'h1ff;
			16'h1f88: y = 16'h1ff;
			16'h1f89: y = 16'h1ff;
			16'h1f8a: y = 16'h1ff;
			16'h1f8b: y = 16'h1ff;
			16'h1f8c: y = 16'h1ff;
			16'h1f8d: y = 16'h1ff;
			16'h1f8e: y = 16'h1ff;
			16'h1f8f: y = 16'h1ff;
			16'h1f90: y = 16'h1ff;
			16'h1f91: y = 16'h1ff;
			16'h1f92: y = 16'h1ff;
			16'h1f93: y = 16'h1ff;
			16'h1f94: y = 16'h1ff;
			16'h1f95: y = 16'h1ff;
			16'h1f96: y = 16'h1ff;
			16'h1f97: y = 16'h1ff;
			16'h1f98: y = 16'h1ff;
			16'h1f99: y = 16'h1ff;
			16'h1f9a: y = 16'h1ff;
			16'h1f9b: y = 16'h1ff;
			16'h1f9c: y = 16'h1ff;
			16'h1f9d: y = 16'h1ff;
			16'h1f9e: y = 16'h1ff;
			16'h1f9f: y = 16'h1ff;
			16'h1fa0: y = 16'h1ff;
			16'h1fa1: y = 16'h1ff;
			16'h1fa2: y = 16'h1ff;
			16'h1fa3: y = 16'h1ff;
			16'h1fa4: y = 16'h1ff;
			16'h1fa5: y = 16'h1ff;
			16'h1fa6: y = 16'h1ff;
			16'h1fa7: y = 16'h1ff;
			16'h1fa8: y = 16'h1ff;
			16'h1fa9: y = 16'h1ff;
			16'h1faa: y = 16'h1ff;
			16'h1fab: y = 16'h1ff;
			16'h1fac: y = 16'h1ff;
			16'h1fad: y = 16'h1ff;
			16'h1fae: y = 16'h1ff;
			16'h1faf: y = 16'h1ff;
			16'h1fb0: y = 16'h1ff;
			16'h1fb1: y = 16'h1ff;
			16'h1fb2: y = 16'h1ff;
			16'h1fb3: y = 16'h1ff;
			16'h1fb4: y = 16'h1ff;
			16'h1fb5: y = 16'h1ff;
			16'h1fb6: y = 16'h1ff;
			16'h1fb7: y = 16'h1ff;
			16'h1fb8: y = 16'h1ff;
			16'h1fb9: y = 16'h1ff;
			16'h1fba: y = 16'h1ff;
			16'h1fbb: y = 16'h1ff;
			16'h1fbc: y = 16'h1ff;
			16'h1fbd: y = 16'h1ff;
			16'h1fbe: y = 16'h1ff;
			16'h1fbf: y = 16'h1ff;
			16'h1fc0: y = 16'h1ff;
			16'h1fc1: y = 16'h1ff;
			16'h1fc2: y = 16'h1ff;
			16'h1fc3: y = 16'h1ff;
			16'h1fc4: y = 16'h1ff;
			16'h1fc5: y = 16'h1ff;
			16'h1fc6: y = 16'h1ff;
			16'h1fc7: y = 16'h1ff;
			16'h1fc8: y = 16'h1ff;
			16'h1fc9: y = 16'h1ff;
			16'h1fca: y = 16'h1ff;
			16'h1fcb: y = 16'h1ff;
			16'h1fcc: y = 16'h1ff;
			16'h1fcd: y = 16'h1ff;
			16'h1fce: y = 16'h1ff;
			16'h1fcf: y = 16'h1ff;
			16'h1fd0: y = 16'h1ff;
			16'h1fd1: y = 16'h1ff;
			16'h1fd2: y = 16'h1ff;
			16'h1fd3: y = 16'h1ff;
			16'h1fd4: y = 16'h1ff;
			16'h1fd5: y = 16'h1ff;
			16'h1fd6: y = 16'h1ff;
			16'h1fd7: y = 16'h1ff;
			16'h1fd8: y = 16'h1ff;
			16'h1fd9: y = 16'h1ff;
			16'h1fda: y = 16'h1ff;
			16'h1fdb: y = 16'h1ff;
			16'h1fdc: y = 16'h1ff;
			16'h1fdd: y = 16'h1ff;
			16'h1fde: y = 16'h1ff;
			16'h1fdf: y = 16'h1ff;
			16'h1fe0: y = 16'h1ff;
			16'h1fe1: y = 16'h1ff;
			16'h1fe2: y = 16'h1ff;
			16'h1fe3: y = 16'h1ff;
			16'h1fe4: y = 16'h1ff;
			16'h1fe5: y = 16'h1ff;
			16'h1fe6: y = 16'h1ff;
			16'h1fe7: y = 16'h1ff;
			16'h1fe8: y = 16'h1ff;
			16'h1fe9: y = 16'h1ff;
			16'h1fea: y = 16'h1ff;
			16'h1feb: y = 16'h1ff;
			16'h1fec: y = 16'h1ff;
			16'h1fed: y = 16'h1ff;
			16'h1fee: y = 16'h1ff;
			16'h1fef: y = 16'h1ff;
			16'h1ff0: y = 16'h1ff;
			16'h1ff1: y = 16'h1ff;
			16'h1ff2: y = 16'h1ff;
			16'h1ff3: y = 16'h1ff;
			16'h1ff4: y = 16'h1ff;
			16'h1ff5: y = 16'h1ff;
			16'h1ff6: y = 16'h1ff;
			16'h1ff7: y = 16'h1ff;
			16'h1ff8: y = 16'h1ff;
			16'h1ff9: y = 16'h1ff;
			16'h1ffa: y = 16'h1ff;
			16'h1ffb: y = 16'h1ff;
			16'h1ffc: y = 16'h1ff;
			16'h1ffd: y = 16'h1ff;
			16'h1ffe: y = 16'h1ff;
			16'h1fff: y = 16'h1ff;
			16'h2000: y = 16'h1ff;
			16'h2001: y = 16'h1ff;
			16'h2002: y = 16'h1ff;
			16'h2003: y = 16'h1ff;
			16'h2004: y = 16'h1ff;
			16'h2005: y = 16'h1ff;
			16'h2006: y = 16'h1ff;
			16'h2007: y = 16'h1ff;
			16'h2008: y = 16'h1ff;
			16'h2009: y = 16'h1ff;
			16'h200a: y = 16'h1ff;
			16'h200b: y = 16'h1ff;
			16'h200c: y = 16'h1ff;
			16'h200d: y = 16'h1ff;
			16'h200e: y = 16'h1ff;
			16'h200f: y = 16'h1ff;
			16'h2010: y = 16'h1ff;
			16'h2011: y = 16'h1ff;
			16'h2012: y = 16'h1ff;
			16'h2013: y = 16'h1ff;
			16'h2014: y = 16'h1ff;
			16'h2015: y = 16'h1ff;
			16'h2016: y = 16'h1ff;
			16'h2017: y = 16'h1ff;
			16'h2018: y = 16'h1ff;
			16'h2019: y = 16'h1ff;
			16'h201a: y = 16'h1ff;
			16'h201b: y = 16'h1ff;
			16'h201c: y = 16'h1ff;
			16'h201d: y = 16'h1ff;
			16'h201e: y = 16'h1ff;
			16'h201f: y = 16'h1ff;
			16'h2020: y = 16'h1ff;
			16'h2021: y = 16'h1ff;
			16'h2022: y = 16'h1ff;
			16'h2023: y = 16'h1ff;
			16'h2024: y = 16'h1ff;
			16'h2025: y = 16'h1ff;
			16'h2026: y = 16'h1ff;
			16'h2027: y = 16'h1ff;
			16'h2028: y = 16'h1ff;
			16'h2029: y = 16'h1ff;
			16'h202a: y = 16'h1ff;
			16'h202b: y = 16'h1ff;
			16'h202c: y = 16'h1ff;
			16'h202d: y = 16'h1ff;
			16'h202e: y = 16'h1ff;
			16'h202f: y = 16'h1ff;
			16'h2030: y = 16'h1ff;
			16'h2031: y = 16'h1ff;
			16'h2032: y = 16'h1ff;
			16'h2033: y = 16'h1ff;
			16'h2034: y = 16'h1ff;
			16'h2035: y = 16'h1ff;
			16'h2036: y = 16'h1ff;
			16'h2037: y = 16'h1ff;
			16'h2038: y = 16'h1ff;
			16'h2039: y = 16'h1ff;
			16'h203a: y = 16'h1ff;
			16'h203b: y = 16'h1ff;
			16'h203c: y = 16'h1ff;
			16'h203d: y = 16'h1ff;
			16'h203e: y = 16'h1ff;
			16'h203f: y = 16'h1ff;
			16'h2040: y = 16'h1ff;
			16'h2041: y = 16'h1ff;
			16'h2042: y = 16'h1ff;
			16'h2043: y = 16'h1ff;
			16'h2044: y = 16'h1ff;
			16'h2045: y = 16'h1ff;
			16'h2046: y = 16'h1ff;
			16'h2047: y = 16'h1ff;
			16'h2048: y = 16'h1ff;
			16'h2049: y = 16'h1ff;
			16'h204a: y = 16'h1ff;
			16'h204b: y = 16'h1ff;
			16'h204c: y = 16'h1ff;
			16'h204d: y = 16'h1ff;
			16'h204e: y = 16'h1ff;
			16'h204f: y = 16'h1ff;
			16'h2050: y = 16'h1ff;
			16'h2051: y = 16'h1ff;
			16'h2052: y = 16'h1ff;
			16'h2053: y = 16'h1ff;
			16'h2054: y = 16'h1ff;
			16'h2055: y = 16'h1ff;
			16'h2056: y = 16'h1ff;
			16'h2057: y = 16'h1ff;
			16'h2058: y = 16'h1ff;
			16'h2059: y = 16'h1ff;
			16'h205a: y = 16'h1ff;
			16'h205b: y = 16'h1ff;
			16'h205c: y = 16'h1ff;
			16'h205d: y = 16'h1ff;
			16'h205e: y = 16'h1ff;
			16'h205f: y = 16'h1ff;
			16'h2060: y = 16'h1ff;
			16'h2061: y = 16'h1ff;
			16'h2062: y = 16'h1ff;
			16'h2063: y = 16'h1ff;
			16'h2064: y = 16'h1ff;
			16'h2065: y = 16'h1ff;
			16'h2066: y = 16'h1ff;
			16'h2067: y = 16'h1ff;
			16'h2068: y = 16'h1ff;
			16'h2069: y = 16'h1ff;
			16'h206a: y = 16'h1ff;
			16'h206b: y = 16'h1ff;
			16'h206c: y = 16'h1ff;
			16'h206d: y = 16'h1ff;
			16'h206e: y = 16'h1ff;
			16'h206f: y = 16'h1ff;
			16'h2070: y = 16'h1ff;
			16'h2071: y = 16'h1ff;
			16'h2072: y = 16'h1ff;
			16'h2073: y = 16'h1ff;
			16'h2074: y = 16'h1ff;
			16'h2075: y = 16'h1ff;
			16'h2076: y = 16'h1ff;
			16'h2077: y = 16'h1ff;
			16'h2078: y = 16'h1ff;
			16'h2079: y = 16'h1ff;
			16'h207a: y = 16'h1ff;
			16'h207b: y = 16'h1ff;
			16'h207c: y = 16'h1ff;
			16'h207d: y = 16'h1ff;
			16'h207e: y = 16'h1ff;
			16'h207f: y = 16'h1ff;
			16'h2080: y = 16'h1ff;
			16'h2081: y = 16'h1ff;
			16'h2082: y = 16'h1ff;
			16'h2083: y = 16'h1ff;
			16'h2084: y = 16'h1ff;
			16'h2085: y = 16'h1ff;
			16'h2086: y = 16'h1ff;
			16'h2087: y = 16'h1ff;
			16'h2088: y = 16'h1ff;
			16'h2089: y = 16'h1ff;
			16'h208a: y = 16'h1ff;
			16'h208b: y = 16'h1ff;
			16'h208c: y = 16'h1ff;
			16'h208d: y = 16'h1ff;
			16'h208e: y = 16'h1ff;
			16'h208f: y = 16'h1ff;
			16'h2090: y = 16'h1ff;
			16'h2091: y = 16'h1ff;
			16'h2092: y = 16'h1ff;
			16'h2093: y = 16'h1ff;
			16'h2094: y = 16'h1ff;
			16'h2095: y = 16'h1ff;
			16'h2096: y = 16'h1ff;
			16'h2097: y = 16'h1ff;
			16'h2098: y = 16'h1ff;
			16'h2099: y = 16'h1ff;
			16'h209a: y = 16'h1ff;
			16'h209b: y = 16'h1ff;
			16'h209c: y = 16'h1ff;
			16'h209d: y = 16'h1ff;
			16'h209e: y = 16'h1ff;
			16'h209f: y = 16'h1ff;
			16'h20a0: y = 16'h1ff;
			16'h20a1: y = 16'h1ff;
			16'h20a2: y = 16'h1ff;
			16'h20a3: y = 16'h1ff;
			16'h20a4: y = 16'h1ff;
			16'h20a5: y = 16'h1ff;
			16'h20a6: y = 16'h1ff;
			16'h20a7: y = 16'h1ff;
			16'h20a8: y = 16'h1ff;
			16'h20a9: y = 16'h1ff;
			16'h20aa: y = 16'h1ff;
			16'h20ab: y = 16'h1ff;
			16'h20ac: y = 16'h1ff;
			16'h20ad: y = 16'h1ff;
			16'h20ae: y = 16'h1ff;
			16'h20af: y = 16'h1ff;
			16'h20b0: y = 16'h1ff;
			16'h20b1: y = 16'h1ff;
			16'h20b2: y = 16'h1ff;
			16'h20b3: y = 16'h1ff;
			16'h20b4: y = 16'h1ff;
			16'h20b5: y = 16'h1ff;
			16'h20b6: y = 16'h1ff;
			16'h20b7: y = 16'h1ff;
			16'h20b8: y = 16'h1ff;
			16'h20b9: y = 16'h1ff;
			16'h20ba: y = 16'h1ff;
			16'h20bb: y = 16'h1ff;
			16'h20bc: y = 16'h1ff;
			16'h20bd: y = 16'h1ff;
			16'h20be: y = 16'h1ff;
			16'h20bf: y = 16'h1ff;
			16'h20c0: y = 16'h1ff;
			16'h20c1: y = 16'h1ff;
			16'h20c2: y = 16'h1ff;
			16'h20c3: y = 16'h1ff;
			16'h20c4: y = 16'h1ff;
			16'h20c5: y = 16'h1ff;
			16'h20c6: y = 16'h1ff;
			16'h20c7: y = 16'h1ff;
			16'h20c8: y = 16'h1ff;
			16'h20c9: y = 16'h1ff;
			16'h20ca: y = 16'h1ff;
			16'h20cb: y = 16'h1ff;
			16'h20cc: y = 16'h1ff;
			16'h20cd: y = 16'h1ff;
			16'h20ce: y = 16'h1ff;
			16'h20cf: y = 16'h1ff;
			16'h20d0: y = 16'h1ff;
			16'h20d1: y = 16'h1ff;
			16'h20d2: y = 16'h1ff;
			16'h20d3: y = 16'h1ff;
			16'h20d4: y = 16'h1ff;
			16'h20d5: y = 16'h1ff;
			16'h20d6: y = 16'h1ff;
			16'h20d7: y = 16'h1ff;
			16'h20d8: y = 16'h1ff;
			16'h20d9: y = 16'h1ff;
			16'h20da: y = 16'h1ff;
			16'h20db: y = 16'h1ff;
			16'h20dc: y = 16'h1ff;
			16'h20dd: y = 16'h1ff;
			16'h20de: y = 16'h1ff;
			16'h20df: y = 16'h1ff;
			16'h20e0: y = 16'h1ff;
			16'h20e1: y = 16'h1ff;
			16'h20e2: y = 16'h1ff;
			16'h20e3: y = 16'h1ff;
			16'h20e4: y = 16'h1ff;
			16'h20e5: y = 16'h1ff;
			16'h20e6: y = 16'h1ff;
			16'h20e7: y = 16'h1ff;
			16'h20e8: y = 16'h1ff;
			16'h20e9: y = 16'h1ff;
			16'h20ea: y = 16'h1ff;
			16'h20eb: y = 16'h1ff;
			16'h20ec: y = 16'h1ff;
			16'h20ed: y = 16'h1ff;
			16'h20ee: y = 16'h1ff;
			16'h20ef: y = 16'h1ff;
			16'h20f0: y = 16'h1ff;
			16'h20f1: y = 16'h1ff;
			16'h20f2: y = 16'h1ff;
			16'h20f3: y = 16'h1ff;
			16'h20f4: y = 16'h1ff;
			16'h20f5: y = 16'h1ff;
			16'h20f6: y = 16'h1ff;
			16'h20f7: y = 16'h1ff;
			16'h20f8: y = 16'h1ff;
			16'h20f9: y = 16'h1ff;
			16'h20fa: y = 16'h1ff;
			16'h20fb: y = 16'h1ff;
			16'h20fc: y = 16'h1ff;
			16'h20fd: y = 16'h1ff;
			16'h20fe: y = 16'h1ff;
			16'h20ff: y = 16'h1ff;
			16'h2100: y = 16'h1ff;
			16'h2101: y = 16'h1ff;
			16'h2102: y = 16'h1ff;
			16'h2103: y = 16'h1ff;
			16'h2104: y = 16'h1ff;
			16'h2105: y = 16'h1ff;
			16'h2106: y = 16'h1ff;
			16'h2107: y = 16'h1ff;
			16'h2108: y = 16'h1ff;
			16'h2109: y = 16'h1ff;
			16'h210a: y = 16'h1ff;
			16'h210b: y = 16'h1ff;
			16'h210c: y = 16'h1ff;
			16'h210d: y = 16'h1ff;
			16'h210e: y = 16'h1ff;
			16'h210f: y = 16'h1ff;
			16'h2110: y = 16'h1ff;
			16'h2111: y = 16'h1ff;
			16'h2112: y = 16'h1ff;
			16'h2113: y = 16'h1ff;
			16'h2114: y = 16'h1ff;
			16'h2115: y = 16'h1ff;
			16'h2116: y = 16'h1ff;
			16'h2117: y = 16'h1ff;
			16'h2118: y = 16'h1ff;
			16'h2119: y = 16'h1ff;
			16'h211a: y = 16'h1ff;
			16'h211b: y = 16'h1ff;
			16'h211c: y = 16'h1ff;
			16'h211d: y = 16'h1ff;
			16'h211e: y = 16'h1ff;
			16'h211f: y = 16'h1ff;
			16'h2120: y = 16'h1ff;
			16'h2121: y = 16'h1ff;
			16'h2122: y = 16'h1ff;
			16'h2123: y = 16'h1ff;
			16'h2124: y = 16'h1ff;
			16'h2125: y = 16'h1ff;
			16'h2126: y = 16'h1ff;
			16'h2127: y = 16'h1ff;
			16'h2128: y = 16'h1ff;
			16'h2129: y = 16'h1ff;
			16'h212a: y = 16'h1ff;
			16'h212b: y = 16'h1ff;
			16'h212c: y = 16'h1ff;
			16'h212d: y = 16'h1ff;
			16'h212e: y = 16'h1ff;
			16'h212f: y = 16'h1ff;
			16'h2130: y = 16'h1ff;
			16'h2131: y = 16'h1ff;
			16'h2132: y = 16'h1ff;
			16'h2133: y = 16'h1ff;
			16'h2134: y = 16'h1ff;
			16'h2135: y = 16'h1ff;
			16'h2136: y = 16'h1ff;
			16'h2137: y = 16'h1ff;
			16'h2138: y = 16'h1ff;
			16'h2139: y = 16'h1ff;
			16'h213a: y = 16'h1ff;
			16'h213b: y = 16'h1ff;
			16'h213c: y = 16'h1ff;
			16'h213d: y = 16'h1ff;
			16'h213e: y = 16'h1ff;
			16'h213f: y = 16'h1ff;
			16'h2140: y = 16'h1ff;
			16'h2141: y = 16'h1ff;
			16'h2142: y = 16'h1ff;
			16'h2143: y = 16'h1ff;
			16'h2144: y = 16'h1ff;
			16'h2145: y = 16'h1ff;
			16'h2146: y = 16'h1ff;
			16'h2147: y = 16'h1ff;
			16'h2148: y = 16'h1ff;
			16'h2149: y = 16'h1ff;
			16'h214a: y = 16'h1ff;
			16'h214b: y = 16'h1ff;
			16'h214c: y = 16'h1ff;
			16'h214d: y = 16'h1ff;
			16'h214e: y = 16'h1ff;
			16'h214f: y = 16'h1ff;
			16'h2150: y = 16'h1ff;
			16'h2151: y = 16'h1ff;
			16'h2152: y = 16'h1ff;
			16'h2153: y = 16'h1ff;
			16'h2154: y = 16'h1ff;
			16'h2155: y = 16'h1ff;
			16'h2156: y = 16'h1ff;
			16'h2157: y = 16'h1ff;
			16'h2158: y = 16'h1ff;
			16'h2159: y = 16'h1ff;
			16'h215a: y = 16'h1ff;
			16'h215b: y = 16'h1ff;
			16'h215c: y = 16'h1ff;
			16'h215d: y = 16'h1ff;
			16'h215e: y = 16'h1ff;
			16'h215f: y = 16'h1ff;
			16'h2160: y = 16'h1ff;
			16'h2161: y = 16'h1ff;
			16'h2162: y = 16'h1ff;
			16'h2163: y = 16'h1ff;
			16'h2164: y = 16'h1ff;
			16'h2165: y = 16'h1ff;
			16'h2166: y = 16'h1ff;
			16'h2167: y = 16'h1ff;
			16'h2168: y = 16'h1ff;
			16'h2169: y = 16'h1ff;
			16'h216a: y = 16'h1ff;
			16'h216b: y = 16'h1ff;
			16'h216c: y = 16'h1ff;
			16'h216d: y = 16'h1ff;
			16'h216e: y = 16'h1ff;
			16'h216f: y = 16'h1ff;
			16'h2170: y = 16'h1ff;
			16'h2171: y = 16'h1ff;
			16'h2172: y = 16'h1ff;
			16'h2173: y = 16'h1ff;
			16'h2174: y = 16'h1ff;
			16'h2175: y = 16'h1ff;
			16'h2176: y = 16'h1ff;
			16'h2177: y = 16'h1ff;
			16'h2178: y = 16'h1ff;
			16'h2179: y = 16'h1ff;
			16'h217a: y = 16'h1ff;
			16'h217b: y = 16'h1ff;
			16'h217c: y = 16'h1ff;
			16'h217d: y = 16'h1ff;
			16'h217e: y = 16'h1ff;
			16'h217f: y = 16'h1ff;
			16'h2180: y = 16'h1ff;
			16'h2181: y = 16'h1ff;
			16'h2182: y = 16'h1ff;
			16'h2183: y = 16'h1ff;
			16'h2184: y = 16'h1ff;
			16'h2185: y = 16'h1ff;
			16'h2186: y = 16'h1ff;
			16'h2187: y = 16'h1ff;
			16'h2188: y = 16'h1ff;
			16'h2189: y = 16'h1ff;
			16'h218a: y = 16'h1ff;
			16'h218b: y = 16'h1ff;
			16'h218c: y = 16'h1ff;
			16'h218d: y = 16'h1ff;
			16'h218e: y = 16'h1ff;
			16'h218f: y = 16'h1ff;
			16'h2190: y = 16'h1ff;
			16'h2191: y = 16'h1ff;
			16'h2192: y = 16'h1ff;
			16'h2193: y = 16'h1ff;
			16'h2194: y = 16'h1ff;
			16'h2195: y = 16'h1ff;
			16'h2196: y = 16'h1ff;
			16'h2197: y = 16'h1ff;
			16'h2198: y = 16'h1ff;
			16'h2199: y = 16'h1ff;
			16'h219a: y = 16'h1ff;
			16'h219b: y = 16'h1ff;
			16'h219c: y = 16'h1ff;
			16'h219d: y = 16'h1ff;
			16'h219e: y = 16'h1ff;
			16'h219f: y = 16'h1ff;
			16'h21a0: y = 16'h1ff;
			16'h21a1: y = 16'h1ff;
			16'h21a2: y = 16'h1ff;
			16'h21a3: y = 16'h1ff;
			16'h21a4: y = 16'h1ff;
			16'h21a5: y = 16'h1ff;
			16'h21a6: y = 16'h1ff;
			16'h21a7: y = 16'h1ff;
			16'h21a8: y = 16'h1ff;
			16'h21a9: y = 16'h1ff;
			16'h21aa: y = 16'h1ff;
			16'h21ab: y = 16'h1ff;
			16'h21ac: y = 16'h1ff;
			16'h21ad: y = 16'h1ff;
			16'h21ae: y = 16'h1ff;
			16'h21af: y = 16'h1ff;
			16'h21b0: y = 16'h1ff;
			16'h21b1: y = 16'h1ff;
			16'h21b2: y = 16'h1ff;
			16'h21b3: y = 16'h1ff;
			16'h21b4: y = 16'h1ff;
			16'h21b5: y = 16'h1ff;
			16'h21b6: y = 16'h1ff;
			16'h21b7: y = 16'h1ff;
			16'h21b8: y = 16'h1ff;
			16'h21b9: y = 16'h1ff;
			16'h21ba: y = 16'h1ff;
			16'h21bb: y = 16'h1ff;
			16'h21bc: y = 16'h1ff;
			16'h21bd: y = 16'h1ff;
			16'h21be: y = 16'h1ff;
			16'h21bf: y = 16'h1ff;
			16'h21c0: y = 16'h1ff;
			16'h21c1: y = 16'h1ff;
			16'h21c2: y = 16'h1ff;
			16'h21c3: y = 16'h1ff;
			16'h21c4: y = 16'h1ff;
			16'h21c5: y = 16'h1ff;
			16'h21c6: y = 16'h1ff;
			16'h21c7: y = 16'h1ff;
			16'h21c8: y = 16'h1ff;
			16'h21c9: y = 16'h1ff;
			16'h21ca: y = 16'h1ff;
			16'h21cb: y = 16'h1ff;
			16'h21cc: y = 16'h1ff;
			16'h21cd: y = 16'h1ff;
			16'h21ce: y = 16'h1ff;
			16'h21cf: y = 16'h1ff;
			16'h21d0: y = 16'h1ff;
			16'h21d1: y = 16'h1ff;
			16'h21d2: y = 16'h1ff;
			16'h21d3: y = 16'h1ff;
			16'h21d4: y = 16'h1ff;
			16'h21d5: y = 16'h1ff;
			16'h21d6: y = 16'h1ff;
			16'h21d7: y = 16'h1ff;
			16'h21d8: y = 16'h1ff;
			16'h21d9: y = 16'h1ff;
			16'h21da: y = 16'h1ff;
			16'h21db: y = 16'h1ff;
			16'h21dc: y = 16'h1ff;
			16'h21dd: y = 16'h1ff;
			16'h21de: y = 16'h1ff;
			16'h21df: y = 16'h1ff;
			16'h21e0: y = 16'h1ff;
			16'h21e1: y = 16'h1ff;
			16'h21e2: y = 16'h1ff;
			16'h21e3: y = 16'h1ff;
			16'h21e4: y = 16'h1ff;
			16'h21e5: y = 16'h1ff;
			16'h21e6: y = 16'h1ff;
			16'h21e7: y = 16'h1ff;
			16'h21e8: y = 16'h1ff;
			16'h21e9: y = 16'h1ff;
			16'h21ea: y = 16'h1ff;
			16'h21eb: y = 16'h1ff;
			16'h21ec: y = 16'h1ff;
			16'h21ed: y = 16'h1ff;
			16'h21ee: y = 16'h1ff;
			16'h21ef: y = 16'h1ff;
			16'h21f0: y = 16'h1ff;
			16'h21f1: y = 16'h1ff;
			16'h21f2: y = 16'h1ff;
			16'h21f3: y = 16'h1ff;
			16'h21f4: y = 16'h1ff;
			16'h21f5: y = 16'h1ff;
			16'h21f6: y = 16'h1ff;
			16'h21f7: y = 16'h1ff;
			16'h21f8: y = 16'h1ff;
			16'h21f9: y = 16'h1ff;
			16'h21fa: y = 16'h1ff;
			16'h21fb: y = 16'h1ff;
			16'h21fc: y = 16'h1ff;
			16'h21fd: y = 16'h1ff;
			16'h21fe: y = 16'h1ff;
			16'h21ff: y = 16'h1ff;
			16'h2200: y = 16'h1ff;
			16'h2201: y = 16'h1ff;
			16'h2202: y = 16'h1ff;
			16'h2203: y = 16'h1ff;
			16'h2204: y = 16'h1ff;
			16'h2205: y = 16'h1ff;
			16'h2206: y = 16'h1ff;
			16'h2207: y = 16'h1ff;
			16'h2208: y = 16'h1ff;
			16'h2209: y = 16'h1ff;
			16'h220a: y = 16'h1ff;
			16'h220b: y = 16'h1ff;
			16'h220c: y = 16'h1ff;
			16'h220d: y = 16'h1ff;
			16'h220e: y = 16'h1ff;
			16'h220f: y = 16'h1ff;
			16'h2210: y = 16'h1ff;
			16'h2211: y = 16'h1ff;
			16'h2212: y = 16'h1ff;
			16'h2213: y = 16'h1ff;
			16'h2214: y = 16'h1ff;
			16'h2215: y = 16'h1ff;
			16'h2216: y = 16'h1ff;
			16'h2217: y = 16'h1ff;
			16'h2218: y = 16'h1ff;
			16'h2219: y = 16'h1ff;
			16'h221a: y = 16'h1ff;
			16'h221b: y = 16'h1ff;
			16'h221c: y = 16'h1ff;
			16'h221d: y = 16'h1ff;
			16'h221e: y = 16'h1ff;
			16'h221f: y = 16'h1ff;
			16'h2220: y = 16'h1ff;
			16'h2221: y = 16'h1ff;
			16'h2222: y = 16'h1ff;
			16'h2223: y = 16'h1ff;
			16'h2224: y = 16'h1ff;
			16'h2225: y = 16'h1ff;
			16'h2226: y = 16'h1ff;
			16'h2227: y = 16'h1ff;
			16'h2228: y = 16'h1ff;
			16'h2229: y = 16'h1ff;
			16'h222a: y = 16'h1ff;
			16'h222b: y = 16'h1ff;
			16'h222c: y = 16'h1ff;
			16'h222d: y = 16'h1ff;
			16'h222e: y = 16'h1ff;
			16'h222f: y = 16'h1ff;
			16'h2230: y = 16'h1ff;
			16'h2231: y = 16'h1ff;
			16'h2232: y = 16'h1ff;
			16'h2233: y = 16'h1ff;
			16'h2234: y = 16'h1ff;
			16'h2235: y = 16'h1ff;
			16'h2236: y = 16'h1ff;
			16'h2237: y = 16'h1ff;
			16'h2238: y = 16'h1ff;
			16'h2239: y = 16'h1ff;
			16'h223a: y = 16'h1ff;
			16'h223b: y = 16'h1ff;
			16'h223c: y = 16'h1ff;
			16'h223d: y = 16'h1ff;
			16'h223e: y = 16'h1ff;
			16'h223f: y = 16'h1ff;
			16'h2240: y = 16'h1ff;
			16'h2241: y = 16'h1ff;
			16'h2242: y = 16'h1ff;
			16'h2243: y = 16'h1ff;
			16'h2244: y = 16'h1ff;
			16'h2245: y = 16'h1ff;
			16'h2246: y = 16'h1ff;
			16'h2247: y = 16'h1ff;
			16'h2248: y = 16'h1ff;
			16'h2249: y = 16'h1ff;
			16'h224a: y = 16'h1ff;
			16'h224b: y = 16'h1ff;
			16'h224c: y = 16'h1ff;
			16'h224d: y = 16'h1ff;
			16'h224e: y = 16'h1ff;
			16'h224f: y = 16'h1ff;
			16'h2250: y = 16'h1ff;
			16'h2251: y = 16'h1ff;
			16'h2252: y = 16'h1ff;
			16'h2253: y = 16'h1ff;
			16'h2254: y = 16'h1ff;
			16'h2255: y = 16'h1ff;
			16'h2256: y = 16'h1ff;
			16'h2257: y = 16'h1ff;
			16'h2258: y = 16'h1ff;
			16'h2259: y = 16'h1ff;
			16'h225a: y = 16'h1ff;
			16'h225b: y = 16'h1ff;
			16'h225c: y = 16'h1ff;
			16'h225d: y = 16'h1ff;
			16'h225e: y = 16'h1ff;
			16'h225f: y = 16'h1ff;
			16'h2260: y = 16'h1ff;
			16'h2261: y = 16'h1ff;
			16'h2262: y = 16'h1ff;
			16'h2263: y = 16'h1ff;
			16'h2264: y = 16'h1ff;
			16'h2265: y = 16'h1ff;
			16'h2266: y = 16'h1ff;
			16'h2267: y = 16'h1ff;
			16'h2268: y = 16'h1ff;
			16'h2269: y = 16'h1ff;
			16'h226a: y = 16'h1ff;
			16'h226b: y = 16'h1ff;
			16'h226c: y = 16'h1ff;
			16'h226d: y = 16'h1ff;
			16'h226e: y = 16'h1ff;
			16'h226f: y = 16'h1ff;
			16'h2270: y = 16'h1ff;
			16'h2271: y = 16'h1ff;
			16'h2272: y = 16'h1ff;
			16'h2273: y = 16'h1ff;
			16'h2274: y = 16'h1ff;
			16'h2275: y = 16'h1ff;
			16'h2276: y = 16'h1ff;
			16'h2277: y = 16'h1ff;
			16'h2278: y = 16'h1ff;
			16'h2279: y = 16'h1ff;
			16'h227a: y = 16'h1ff;
			16'h227b: y = 16'h1ff;
			16'h227c: y = 16'h1ff;
			16'h227d: y = 16'h1ff;
			16'h227e: y = 16'h1ff;
			16'h227f: y = 16'h1ff;
			16'h2280: y = 16'h1ff;
			16'h2281: y = 16'h1ff;
			16'h2282: y = 16'h1ff;
			16'h2283: y = 16'h1ff;
			16'h2284: y = 16'h1ff;
			16'h2285: y = 16'h1ff;
			16'h2286: y = 16'h1ff;
			16'h2287: y = 16'h1ff;
			16'h2288: y = 16'h1ff;
			16'h2289: y = 16'h1ff;
			16'h228a: y = 16'h1ff;
			16'h228b: y = 16'h1ff;
			16'h228c: y = 16'h1ff;
			16'h228d: y = 16'h1ff;
			16'h228e: y = 16'h1ff;
			16'h228f: y = 16'h1ff;
			16'h2290: y = 16'h1ff;
			16'h2291: y = 16'h1ff;
			16'h2292: y = 16'h1ff;
			16'h2293: y = 16'h1ff;
			16'h2294: y = 16'h1ff;
			16'h2295: y = 16'h1ff;
			16'h2296: y = 16'h1ff;
			16'h2297: y = 16'h1ff;
			16'h2298: y = 16'h1ff;
			16'h2299: y = 16'h1ff;
			16'h229a: y = 16'h1ff;
			16'h229b: y = 16'h1ff;
			16'h229c: y = 16'h1ff;
			16'h229d: y = 16'h1ff;
			16'h229e: y = 16'h1ff;
			16'h229f: y = 16'h1ff;
			16'h22a0: y = 16'h1ff;
			16'h22a1: y = 16'h1ff;
			16'h22a2: y = 16'h1ff;
			16'h22a3: y = 16'h1ff;
			16'h22a4: y = 16'h1ff;
			16'h22a5: y = 16'h1ff;
			16'h22a6: y = 16'h1ff;
			16'h22a7: y = 16'h1ff;
			16'h22a8: y = 16'h1ff;
			16'h22a9: y = 16'h1ff;
			16'h22aa: y = 16'h1ff;
			16'h22ab: y = 16'h1ff;
			16'h22ac: y = 16'h1ff;
			16'h22ad: y = 16'h1ff;
			16'h22ae: y = 16'h1ff;
			16'h22af: y = 16'h1ff;
			16'h22b0: y = 16'h1ff;
			16'h22b1: y = 16'h1ff;
			16'h22b2: y = 16'h1ff;
			16'h22b3: y = 16'h1ff;
			16'h22b4: y = 16'h1ff;
			16'h22b5: y = 16'h1ff;
			16'h22b6: y = 16'h1ff;
			16'h22b7: y = 16'h1ff;
			16'h22b8: y = 16'h1ff;
			16'h22b9: y = 16'h1ff;
			16'h22ba: y = 16'h1ff;
			16'h22bb: y = 16'h1ff;
			16'h22bc: y = 16'h1ff;
			16'h22bd: y = 16'h1ff;
			16'h22be: y = 16'h1ff;
			16'h22bf: y = 16'h1ff;
			16'h22c0: y = 16'h1ff;
			16'h22c1: y = 16'h1ff;
			16'h22c2: y = 16'h1ff;
			16'h22c3: y = 16'h1ff;
			16'h22c4: y = 16'h1ff;
			16'h22c5: y = 16'h1ff;
			16'h22c6: y = 16'h1ff;
			16'h22c7: y = 16'h1ff;
			16'h22c8: y = 16'h1ff;
			16'h22c9: y = 16'h1ff;
			16'h22ca: y = 16'h1ff;
			16'h22cb: y = 16'h1ff;
			16'h22cc: y = 16'h1ff;
			16'h22cd: y = 16'h1ff;
			16'h22ce: y = 16'h1ff;
			16'h22cf: y = 16'h1ff;
			16'h22d0: y = 16'h1ff;
			16'h22d1: y = 16'h1ff;
			16'h22d2: y = 16'h1ff;
			16'h22d3: y = 16'h1ff;
			16'h22d4: y = 16'h1ff;
			16'h22d5: y = 16'h1ff;
			16'h22d6: y = 16'h1ff;
			16'h22d7: y = 16'h1ff;
			16'h22d8: y = 16'h1ff;
			16'h22d9: y = 16'h1ff;
			16'h22da: y = 16'h1ff;
			16'h22db: y = 16'h1ff;
			16'h22dc: y = 16'h1ff;
			16'h22dd: y = 16'h1ff;
			16'h22de: y = 16'h1ff;
			16'h22df: y = 16'h1ff;
			16'h22e0: y = 16'h1ff;
			16'h22e1: y = 16'h1ff;
			16'h22e2: y = 16'h1ff;
			16'h22e3: y = 16'h1ff;
			16'h22e4: y = 16'h1ff;
			16'h22e5: y = 16'h1ff;
			16'h22e6: y = 16'h1ff;
			16'h22e7: y = 16'h1ff;
			16'h22e8: y = 16'h1ff;
			16'h22e9: y = 16'h1ff;
			16'h22ea: y = 16'h1ff;
			16'h22eb: y = 16'h1ff;
			16'h22ec: y = 16'h1ff;
			16'h22ed: y = 16'h1ff;
			16'h22ee: y = 16'h1ff;
			16'h22ef: y = 16'h1ff;
			16'h22f0: y = 16'h1ff;
			16'h22f1: y = 16'h1ff;
			16'h22f2: y = 16'h1ff;
			16'h22f3: y = 16'h1ff;
			16'h22f4: y = 16'h1ff;
			16'h22f5: y = 16'h1ff;
			16'h22f6: y = 16'h1ff;
			16'h22f7: y = 16'h1ff;
			16'h22f8: y = 16'h1ff;
			16'h22f9: y = 16'h1ff;
			16'h22fa: y = 16'h1ff;
			16'h22fb: y = 16'h1ff;
			16'h22fc: y = 16'h1ff;
			16'h22fd: y = 16'h1ff;
			16'h22fe: y = 16'h1ff;
			16'h22ff: y = 16'h1ff;
			16'h2300: y = 16'h1ff;
			16'h2301: y = 16'h1ff;
			16'h2302: y = 16'h1ff;
			16'h2303: y = 16'h1ff;
			16'h2304: y = 16'h1ff;
			16'h2305: y = 16'h1ff;
			16'h2306: y = 16'h1ff;
			16'h2307: y = 16'h1ff;
			16'h2308: y = 16'h1ff;
			16'h2309: y = 16'h1ff;
			16'h230a: y = 16'h1ff;
			16'h230b: y = 16'h1ff;
			16'h230c: y = 16'h1ff;
			16'h230d: y = 16'h1ff;
			16'h230e: y = 16'h1ff;
			16'h230f: y = 16'h1ff;
			16'h2310: y = 16'h1ff;
			16'h2311: y = 16'h1ff;
			16'h2312: y = 16'h1ff;
			16'h2313: y = 16'h1ff;
			16'h2314: y = 16'h1ff;
			16'h2315: y = 16'h1ff;
			16'h2316: y = 16'h1ff;
			16'h2317: y = 16'h1ff;
			16'h2318: y = 16'h1ff;
			16'h2319: y = 16'h1ff;
			16'h231a: y = 16'h1ff;
			16'h231b: y = 16'h1ff;
			16'h231c: y = 16'h1ff;
			16'h231d: y = 16'h1ff;
			16'h231e: y = 16'h1ff;
			16'h231f: y = 16'h1ff;
			16'h2320: y = 16'h1ff;
			16'h2321: y = 16'h1ff;
			16'h2322: y = 16'h1ff;
			16'h2323: y = 16'h1ff;
			16'h2324: y = 16'h1ff;
			16'h2325: y = 16'h1ff;
			16'h2326: y = 16'h1ff;
			16'h2327: y = 16'h1ff;
			16'h2328: y = 16'h1ff;
			16'h2329: y = 16'h1ff;
			16'h232a: y = 16'h1ff;
			16'h232b: y = 16'h1ff;
			16'h232c: y = 16'h1ff;
			16'h232d: y = 16'h1ff;
			16'h232e: y = 16'h1ff;
			16'h232f: y = 16'h1ff;
			16'h2330: y = 16'h1ff;
			16'h2331: y = 16'h1ff;
			16'h2332: y = 16'h1ff;
			16'h2333: y = 16'h1ff;
			16'h2334: y = 16'h1ff;
			16'h2335: y = 16'h1ff;
			16'h2336: y = 16'h1ff;
			16'h2337: y = 16'h1ff;
			16'h2338: y = 16'h1ff;
			16'h2339: y = 16'h1ff;
			16'h233a: y = 16'h1ff;
			16'h233b: y = 16'h1ff;
			16'h233c: y = 16'h1ff;
			16'h233d: y = 16'h1ff;
			16'h233e: y = 16'h1ff;
			16'h233f: y = 16'h1ff;
			16'h2340: y = 16'h1ff;
			16'h2341: y = 16'h1ff;
			16'h2342: y = 16'h1ff;
			16'h2343: y = 16'h1ff;
			16'h2344: y = 16'h1ff;
			16'h2345: y = 16'h1ff;
			16'h2346: y = 16'h1ff;
			16'h2347: y = 16'h1ff;
			16'h2348: y = 16'h1ff;
			16'h2349: y = 16'h1ff;
			16'h234a: y = 16'h1ff;
			16'h234b: y = 16'h1ff;
			16'h234c: y = 16'h1ff;
			16'h234d: y = 16'h1ff;
			16'h234e: y = 16'h1ff;
			16'h234f: y = 16'h1ff;
			16'h2350: y = 16'h1ff;
			16'h2351: y = 16'h1ff;
			16'h2352: y = 16'h1ff;
			16'h2353: y = 16'h1ff;
			16'h2354: y = 16'h1ff;
			16'h2355: y = 16'h1ff;
			16'h2356: y = 16'h1ff;
			16'h2357: y = 16'h1ff;
			16'h2358: y = 16'h1ff;
			16'h2359: y = 16'h1ff;
			16'h235a: y = 16'h1ff;
			16'h235b: y = 16'h1ff;
			16'h235c: y = 16'h1ff;
			16'h235d: y = 16'h1ff;
			16'h235e: y = 16'h1ff;
			16'h235f: y = 16'h1ff;
			16'h2360: y = 16'h1ff;
			16'h2361: y = 16'h1ff;
			16'h2362: y = 16'h1ff;
			16'h2363: y = 16'h1ff;
			16'h2364: y = 16'h1ff;
			16'h2365: y = 16'h1ff;
			16'h2366: y = 16'h1ff;
			16'h2367: y = 16'h1ff;
			16'h2368: y = 16'h1ff;
			16'h2369: y = 16'h1ff;
			16'h236a: y = 16'h1ff;
			16'h236b: y = 16'h1ff;
			16'h236c: y = 16'h1ff;
			16'h236d: y = 16'h1ff;
			16'h236e: y = 16'h1ff;
			16'h236f: y = 16'h1ff;
			16'h2370: y = 16'h1ff;
			16'h2371: y = 16'h1ff;
			16'h2372: y = 16'h1ff;
			16'h2373: y = 16'h1ff;
			16'h2374: y = 16'h1ff;
			16'h2375: y = 16'h1ff;
			16'h2376: y = 16'h1ff;
			16'h2377: y = 16'h1ff;
			16'h2378: y = 16'h1ff;
			16'h2379: y = 16'h1ff;
			16'h237a: y = 16'h1ff;
			16'h237b: y = 16'h1ff;
			16'h237c: y = 16'h1ff;
			16'h237d: y = 16'h1ff;
			16'h237e: y = 16'h1ff;
			16'h237f: y = 16'h1ff;
			16'h2380: y = 16'h1ff;
			16'h2381: y = 16'h1ff;
			16'h2382: y = 16'h1ff;
			16'h2383: y = 16'h1ff;
			16'h2384: y = 16'h1ff;
			16'h2385: y = 16'h1ff;
			16'h2386: y = 16'h1ff;
			16'h2387: y = 16'h1ff;
			16'h2388: y = 16'h1ff;
			16'h2389: y = 16'h1ff;
			16'h238a: y = 16'h1ff;
			16'h238b: y = 16'h1ff;
			16'h238c: y = 16'h1ff;
			16'h238d: y = 16'h1ff;
			16'h238e: y = 16'h1ff;
			16'h238f: y = 16'h1ff;
			16'h2390: y = 16'h1ff;
			16'h2391: y = 16'h1ff;
			16'h2392: y = 16'h1ff;
			16'h2393: y = 16'h1ff;
			16'h2394: y = 16'h1ff;
			16'h2395: y = 16'h1ff;
			16'h2396: y = 16'h1ff;
			16'h2397: y = 16'h1ff;
			16'h2398: y = 16'h1ff;
			16'h2399: y = 16'h1ff;
			16'h239a: y = 16'h1ff;
			16'h239b: y = 16'h1ff;
			16'h239c: y = 16'h1ff;
			16'h239d: y = 16'h1ff;
			16'h239e: y = 16'h1ff;
			16'h239f: y = 16'h1ff;
			16'h23a0: y = 16'h1ff;
			16'h23a1: y = 16'h1ff;
			16'h23a2: y = 16'h1ff;
			16'h23a3: y = 16'h1ff;
			16'h23a4: y = 16'h1ff;
			16'h23a5: y = 16'h1ff;
			16'h23a6: y = 16'h1ff;
			16'h23a7: y = 16'h1ff;
			16'h23a8: y = 16'h1ff;
			16'h23a9: y = 16'h1ff;
			16'h23aa: y = 16'h1ff;
			16'h23ab: y = 16'h1ff;
			16'h23ac: y = 16'h1ff;
			16'h23ad: y = 16'h1ff;
			16'h23ae: y = 16'h1ff;
			16'h23af: y = 16'h1ff;
			16'h23b0: y = 16'h1ff;
			16'h23b1: y = 16'h1ff;
			16'h23b2: y = 16'h1ff;
			16'h23b3: y = 16'h1ff;
			16'h23b4: y = 16'h1ff;
			16'h23b5: y = 16'h1ff;
			16'h23b6: y = 16'h1ff;
			16'h23b7: y = 16'h1ff;
			16'h23b8: y = 16'h1ff;
			16'h23b9: y = 16'h1ff;
			16'h23ba: y = 16'h1ff;
			16'h23bb: y = 16'h1ff;
			16'h23bc: y = 16'h1ff;
			16'h23bd: y = 16'h1ff;
			16'h23be: y = 16'h1ff;
			16'h23bf: y = 16'h1ff;
			16'h23c0: y = 16'h1ff;
			16'h23c1: y = 16'h1ff;
			16'h23c2: y = 16'h1ff;
			16'h23c3: y = 16'h1ff;
			16'h23c4: y = 16'h1ff;
			16'h23c5: y = 16'h1ff;
			16'h23c6: y = 16'h1ff;
			16'h23c7: y = 16'h1ff;
			16'h23c8: y = 16'h1ff;
			16'h23c9: y = 16'h1ff;
			16'h23ca: y = 16'h1ff;
			16'h23cb: y = 16'h1ff;
			16'h23cc: y = 16'h1ff;
			16'h23cd: y = 16'h1ff;
			16'h23ce: y = 16'h1ff;
			16'h23cf: y = 16'h1ff;
			16'h23d0: y = 16'h1ff;
			16'h23d1: y = 16'h1ff;
			16'h23d2: y = 16'h1ff;
			16'h23d3: y = 16'h1ff;
			16'h23d4: y = 16'h1ff;
			16'h23d5: y = 16'h1ff;
			16'h23d6: y = 16'h1ff;
			16'h23d7: y = 16'h1ff;
			16'h23d8: y = 16'h1ff;
			16'h23d9: y = 16'h1ff;
			16'h23da: y = 16'h1ff;
			16'h23db: y = 16'h1ff;
			16'h23dc: y = 16'h1ff;
			16'h23dd: y = 16'h1ff;
			16'h23de: y = 16'h1ff;
			16'h23df: y = 16'h1ff;
			16'h23e0: y = 16'h1ff;
			16'h23e1: y = 16'h1ff;
			16'h23e2: y = 16'h1ff;
			16'h23e3: y = 16'h1ff;
			16'h23e4: y = 16'h1ff;
			16'h23e5: y = 16'h1ff;
			16'h23e6: y = 16'h1ff;
			16'h23e7: y = 16'h1ff;
			16'h23e8: y = 16'h1ff;
			16'h23e9: y = 16'h1ff;
			16'h23ea: y = 16'h1ff;
			16'h23eb: y = 16'h1ff;
			16'h23ec: y = 16'h1ff;
			16'h23ed: y = 16'h1ff;
			16'h23ee: y = 16'h1ff;
			16'h23ef: y = 16'h1ff;
			16'h23f0: y = 16'h1ff;
			16'h23f1: y = 16'h1ff;
			16'h23f2: y = 16'h1ff;
			16'h23f3: y = 16'h1ff;
			16'h23f4: y = 16'h1ff;
			16'h23f5: y = 16'h1ff;
			16'h23f6: y = 16'h1ff;
			16'h23f7: y = 16'h1ff;
			16'h23f8: y = 16'h1ff;
			16'h23f9: y = 16'h1ff;
			16'h23fa: y = 16'h1ff;
			16'h23fb: y = 16'h1ff;
			16'h23fc: y = 16'h1ff;
			16'h23fd: y = 16'h1ff;
			16'h23fe: y = 16'h1ff;
			16'h23ff: y = 16'h1ff;
			16'h2400: y = 16'h1ff;
			16'h2401: y = 16'h1ff;
			16'h2402: y = 16'h1ff;
			16'h2403: y = 16'h1ff;
			16'h2404: y = 16'h1ff;
			16'h2405: y = 16'h1ff;
			16'h2406: y = 16'h1ff;
			16'h2407: y = 16'h1ff;
			16'h2408: y = 16'h1ff;
			16'h2409: y = 16'h1ff;
			16'h240a: y = 16'h1ff;
			16'h240b: y = 16'h1ff;
			16'h240c: y = 16'h1ff;
			16'h240d: y = 16'h1ff;
			16'h240e: y = 16'h1ff;
			16'h240f: y = 16'h1ff;
			16'h2410: y = 16'h1ff;
			16'h2411: y = 16'h1ff;
			16'h2412: y = 16'h1ff;
			16'h2413: y = 16'h1ff;
			16'h2414: y = 16'h1ff;
			16'h2415: y = 16'h1ff;
			16'h2416: y = 16'h1ff;
			16'h2417: y = 16'h1ff;
			16'h2418: y = 16'h1ff;
			16'h2419: y = 16'h1ff;
			16'h241a: y = 16'h1ff;
			16'h241b: y = 16'h1ff;
			16'h241c: y = 16'h1ff;
			16'h241d: y = 16'h1ff;
			16'h241e: y = 16'h1ff;
			16'h241f: y = 16'h1ff;
			16'h2420: y = 16'h1ff;
			16'h2421: y = 16'h1ff;
			16'h2422: y = 16'h1ff;
			16'h2423: y = 16'h1ff;
			16'h2424: y = 16'h1ff;
			16'h2425: y = 16'h1ff;
			16'h2426: y = 16'h1ff;
			16'h2427: y = 16'h1ff;
			16'h2428: y = 16'h1ff;
			16'h2429: y = 16'h1ff;
			16'h242a: y = 16'h1ff;
			16'h242b: y = 16'h1ff;
			16'h242c: y = 16'h1ff;
			16'h242d: y = 16'h1ff;
			16'h242e: y = 16'h1ff;
			16'h242f: y = 16'h1ff;
			16'h2430: y = 16'h1ff;
			16'h2431: y = 16'h1ff;
			16'h2432: y = 16'h1ff;
			16'h2433: y = 16'h1ff;
			16'h2434: y = 16'h1ff;
			16'h2435: y = 16'h1ff;
			16'h2436: y = 16'h1ff;
			16'h2437: y = 16'h1ff;
			16'h2438: y = 16'h1ff;
			16'h2439: y = 16'h1ff;
			16'h243a: y = 16'h1ff;
			16'h243b: y = 16'h1ff;
			16'h243c: y = 16'h1ff;
			16'h243d: y = 16'h1ff;
			16'h243e: y = 16'h1ff;
			16'h243f: y = 16'h1ff;
			16'h2440: y = 16'h1ff;
			16'h2441: y = 16'h1ff;
			16'h2442: y = 16'h1ff;
			16'h2443: y = 16'h1ff;
			16'h2444: y = 16'h1ff;
			16'h2445: y = 16'h1ff;
			16'h2446: y = 16'h1ff;
			16'h2447: y = 16'h1ff;
			16'h2448: y = 16'h1ff;
			16'h2449: y = 16'h1ff;
			16'h244a: y = 16'h1ff;
			16'h244b: y = 16'h1ff;
			16'h244c: y = 16'h1ff;
			16'h244d: y = 16'h1ff;
			16'h244e: y = 16'h1ff;
			16'h244f: y = 16'h1ff;
			16'h2450: y = 16'h1ff;
			16'h2451: y = 16'h1ff;
			16'h2452: y = 16'h1ff;
			16'h2453: y = 16'h1ff;
			16'h2454: y = 16'h1ff;
			16'h2455: y = 16'h1ff;
			16'h2456: y = 16'h1ff;
			16'h2457: y = 16'h1ff;
			16'h2458: y = 16'h1ff;
			16'h2459: y = 16'h1ff;
			16'h245a: y = 16'h1ff;
			16'h245b: y = 16'h1ff;
			16'h245c: y = 16'h1ff;
			16'h245d: y = 16'h1ff;
			16'h245e: y = 16'h1ff;
			16'h245f: y = 16'h1ff;
			16'h2460: y = 16'h1ff;
			16'h2461: y = 16'h1ff;
			16'h2462: y = 16'h1ff;
			16'h2463: y = 16'h1ff;
			16'h2464: y = 16'h1ff;
			16'h2465: y = 16'h1ff;
			16'h2466: y = 16'h1ff;
			16'h2467: y = 16'h1ff;
			16'h2468: y = 16'h1ff;
			16'h2469: y = 16'h1ff;
			16'h246a: y = 16'h1ff;
			16'h246b: y = 16'h1ff;
			16'h246c: y = 16'h1ff;
			16'h246d: y = 16'h1ff;
			16'h246e: y = 16'h1ff;
			16'h246f: y = 16'h1ff;
			16'h2470: y = 16'h1ff;
			16'h2471: y = 16'h1ff;
			16'h2472: y = 16'h1ff;
			16'h2473: y = 16'h1ff;
			16'h2474: y = 16'h1ff;
			16'h2475: y = 16'h1ff;
			16'h2476: y = 16'h1ff;
			16'h2477: y = 16'h1ff;
			16'h2478: y = 16'h1ff;
			16'h2479: y = 16'h1ff;
			16'h247a: y = 16'h1ff;
			16'h247b: y = 16'h1ff;
			16'h247c: y = 16'h1ff;
			16'h247d: y = 16'h1ff;
			16'h247e: y = 16'h1ff;
			16'h247f: y = 16'h1ff;
			16'h2480: y = 16'h1ff;
			16'h2481: y = 16'h1ff;
			16'h2482: y = 16'h1ff;
			16'h2483: y = 16'h1ff;
			16'h2484: y = 16'h1ff;
			16'h2485: y = 16'h1ff;
			16'h2486: y = 16'h1ff;
			16'h2487: y = 16'h1ff;
			16'h2488: y = 16'h1ff;
			16'h2489: y = 16'h1ff;
			16'h248a: y = 16'h1ff;
			16'h248b: y = 16'h1ff;
			16'h248c: y = 16'h1ff;
			16'h248d: y = 16'h1ff;
			16'h248e: y = 16'h1ff;
			16'h248f: y = 16'h1ff;
			16'h2490: y = 16'h1ff;
			16'h2491: y = 16'h1ff;
			16'h2492: y = 16'h1ff;
			16'h2493: y = 16'h1ff;
			16'h2494: y = 16'h1ff;
			16'h2495: y = 16'h1ff;
			16'h2496: y = 16'h1ff;
			16'h2497: y = 16'h1ff;
			16'h2498: y = 16'h1ff;
			16'h2499: y = 16'h1ff;
			16'h249a: y = 16'h1ff;
			16'h249b: y = 16'h1ff;
			16'h249c: y = 16'h1ff;
			16'h249d: y = 16'h1ff;
			16'h249e: y = 16'h1ff;
			16'h249f: y = 16'h1ff;
			16'h24a0: y = 16'h1ff;
			16'h24a1: y = 16'h1ff;
			16'h24a2: y = 16'h1ff;
			16'h24a3: y = 16'h1ff;
			16'h24a4: y = 16'h1ff;
			16'h24a5: y = 16'h1ff;
			16'h24a6: y = 16'h1ff;
			16'h24a7: y = 16'h1ff;
			16'h24a8: y = 16'h1ff;
			16'h24a9: y = 16'h1ff;
			16'h24aa: y = 16'h1ff;
			16'h24ab: y = 16'h1ff;
			16'h24ac: y = 16'h1ff;
			16'h24ad: y = 16'h1ff;
			16'h24ae: y = 16'h1ff;
			16'h24af: y = 16'h1ff;
			16'h24b0: y = 16'h1ff;
			16'h24b1: y = 16'h1ff;
			16'h24b2: y = 16'h1ff;
			16'h24b3: y = 16'h1ff;
			16'h24b4: y = 16'h1ff;
			16'h24b5: y = 16'h1ff;
			16'h24b6: y = 16'h1ff;
			16'h24b7: y = 16'h1ff;
			16'h24b8: y = 16'h1ff;
			16'h24b9: y = 16'h1ff;
			16'h24ba: y = 16'h1ff;
			16'h24bb: y = 16'h1ff;
			16'h24bc: y = 16'h1ff;
			16'h24bd: y = 16'h1ff;
			16'h24be: y = 16'h1ff;
			16'h24bf: y = 16'h1ff;
			16'h24c0: y = 16'h1ff;
			16'h24c1: y = 16'h1ff;
			16'h24c2: y = 16'h1ff;
			16'h24c3: y = 16'h1ff;
			16'h24c4: y = 16'h1ff;
			16'h24c5: y = 16'h1ff;
			16'h24c6: y = 16'h1ff;
			16'h24c7: y = 16'h1ff;
			16'h24c8: y = 16'h1ff;
			16'h24c9: y = 16'h1ff;
			16'h24ca: y = 16'h1ff;
			16'h24cb: y = 16'h1ff;
			16'h24cc: y = 16'h1ff;
			16'h24cd: y = 16'h1ff;
			16'h24ce: y = 16'h1ff;
			16'h24cf: y = 16'h1ff;
			16'h24d0: y = 16'h1ff;
			16'h24d1: y = 16'h1ff;
			16'h24d2: y = 16'h1ff;
			16'h24d3: y = 16'h1ff;
			16'h24d4: y = 16'h1ff;
			16'h24d5: y = 16'h1ff;
			16'h24d6: y = 16'h1ff;
			16'h24d7: y = 16'h1ff;
			16'h24d8: y = 16'h1ff;
			16'h24d9: y = 16'h1ff;
			16'h24da: y = 16'h1ff;
			16'h24db: y = 16'h1ff;
			16'h24dc: y = 16'h1ff;
			16'h24dd: y = 16'h1ff;
			16'h24de: y = 16'h1ff;
			16'h24df: y = 16'h1ff;
			16'h24e0: y = 16'h1ff;
			16'h24e1: y = 16'h1ff;
			16'h24e2: y = 16'h1ff;
			16'h24e3: y = 16'h1ff;
			16'h24e4: y = 16'h1ff;
			16'h24e5: y = 16'h1ff;
			16'h24e6: y = 16'h1ff;
			16'h24e7: y = 16'h1ff;
			16'h24e8: y = 16'h1ff;
			16'h24e9: y = 16'h1ff;
			16'h24ea: y = 16'h1ff;
			16'h24eb: y = 16'h1ff;
			16'h24ec: y = 16'h1ff;
			16'h24ed: y = 16'h1ff;
			16'h24ee: y = 16'h1ff;
			16'h24ef: y = 16'h1ff;
			16'h24f0: y = 16'h1ff;
			16'h24f1: y = 16'h1ff;
			16'h24f2: y = 16'h1ff;
			16'h24f3: y = 16'h1ff;
			16'h24f4: y = 16'h1ff;
			16'h24f5: y = 16'h1ff;
			16'h24f6: y = 16'h1ff;
			16'h24f7: y = 16'h1ff;
			16'h24f8: y = 16'h1ff;
			16'h24f9: y = 16'h1ff;
			16'h24fa: y = 16'h1ff;
			16'h24fb: y = 16'h1ff;
			16'h24fc: y = 16'h1ff;
			16'h24fd: y = 16'h1ff;
			16'h24fe: y = 16'h1ff;
			16'h24ff: y = 16'h1ff;
			16'h2500: y = 16'h1ff;
			16'h2501: y = 16'h1ff;
			16'h2502: y = 16'h1ff;
			16'h2503: y = 16'h1ff;
			16'h2504: y = 16'h1ff;
			16'h2505: y = 16'h1ff;
			16'h2506: y = 16'h1ff;
			16'h2507: y = 16'h1ff;
			16'h2508: y = 16'h1ff;
			16'h2509: y = 16'h1ff;
			16'h250a: y = 16'h1ff;
			16'h250b: y = 16'h1ff;
			16'h250c: y = 16'h1ff;
			16'h250d: y = 16'h1ff;
			16'h250e: y = 16'h1ff;
			16'h250f: y = 16'h1ff;
			16'h2510: y = 16'h1ff;
			16'h2511: y = 16'h1ff;
			16'h2512: y = 16'h1ff;
			16'h2513: y = 16'h1ff;
			16'h2514: y = 16'h1ff;
			16'h2515: y = 16'h1ff;
			16'h2516: y = 16'h1ff;
			16'h2517: y = 16'h1ff;
			16'h2518: y = 16'h1ff;
			16'h2519: y = 16'h1ff;
			16'h251a: y = 16'h1ff;
			16'h251b: y = 16'h1ff;
			16'h251c: y = 16'h1ff;
			16'h251d: y = 16'h1ff;
			16'h251e: y = 16'h1ff;
			16'h251f: y = 16'h1ff;
			16'h2520: y = 16'h1ff;
			16'h2521: y = 16'h1ff;
			16'h2522: y = 16'h1ff;
			16'h2523: y = 16'h1ff;
			16'h2524: y = 16'h1ff;
			16'h2525: y = 16'h1ff;
			16'h2526: y = 16'h1ff;
			16'h2527: y = 16'h1ff;
			16'h2528: y = 16'h1ff;
			16'h2529: y = 16'h1ff;
			16'h252a: y = 16'h1ff;
			16'h252b: y = 16'h1ff;
			16'h252c: y = 16'h1ff;
			16'h252d: y = 16'h1ff;
			16'h252e: y = 16'h1ff;
			16'h252f: y = 16'h1ff;
			16'h2530: y = 16'h1ff;
			16'h2531: y = 16'h1ff;
			16'h2532: y = 16'h1ff;
			16'h2533: y = 16'h1ff;
			16'h2534: y = 16'h1ff;
			16'h2535: y = 16'h1ff;
			16'h2536: y = 16'h1ff;
			16'h2537: y = 16'h1ff;
			16'h2538: y = 16'h1ff;
			16'h2539: y = 16'h1ff;
			16'h253a: y = 16'h1ff;
			16'h253b: y = 16'h1ff;
			16'h253c: y = 16'h1ff;
			16'h253d: y = 16'h1ff;
			16'h253e: y = 16'h1ff;
			16'h253f: y = 16'h1ff;
			16'h2540: y = 16'h1ff;
			16'h2541: y = 16'h1ff;
			16'h2542: y = 16'h1ff;
			16'h2543: y = 16'h1ff;
			16'h2544: y = 16'h1ff;
			16'h2545: y = 16'h1ff;
			16'h2546: y = 16'h1ff;
			16'h2547: y = 16'h1ff;
			16'h2548: y = 16'h1ff;
			16'h2549: y = 16'h1ff;
			16'h254a: y = 16'h1ff;
			16'h254b: y = 16'h1ff;
			16'h254c: y = 16'h1ff;
			16'h254d: y = 16'h1ff;
			16'h254e: y = 16'h1ff;
			16'h254f: y = 16'h1ff;
			16'h2550: y = 16'h1ff;
			16'h2551: y = 16'h1ff;
			16'h2552: y = 16'h1ff;
			16'h2553: y = 16'h1ff;
			16'h2554: y = 16'h1ff;
			16'h2555: y = 16'h1ff;
			16'h2556: y = 16'h1ff;
			16'h2557: y = 16'h1ff;
			16'h2558: y = 16'h1ff;
			16'h2559: y = 16'h1ff;
			16'h255a: y = 16'h1ff;
			16'h255b: y = 16'h1ff;
			16'h255c: y = 16'h1ff;
			16'h255d: y = 16'h1ff;
			16'h255e: y = 16'h1ff;
			16'h255f: y = 16'h1ff;
			16'h2560: y = 16'h1ff;
			16'h2561: y = 16'h1ff;
			16'h2562: y = 16'h1ff;
			16'h2563: y = 16'h1ff;
			16'h2564: y = 16'h1ff;
			16'h2565: y = 16'h1ff;
			16'h2566: y = 16'h1ff;
			16'h2567: y = 16'h1ff;
			16'h2568: y = 16'h1ff;
			16'h2569: y = 16'h1ff;
			16'h256a: y = 16'h1ff;
			16'h256b: y = 16'h1ff;
			16'h256c: y = 16'h1ff;
			16'h256d: y = 16'h1ff;
			16'h256e: y = 16'h1ff;
			16'h256f: y = 16'h200;
			16'h2570: y = 16'h200;
			16'h2571: y = 16'h200;
			16'h2572: y = 16'h200;
			16'h2573: y = 16'h200;
			16'h2574: y = 16'h200;
			16'h2575: y = 16'h200;
			16'h2576: y = 16'h200;
			16'h2577: y = 16'h200;
			16'h2578: y = 16'h200;
			16'h2579: y = 16'h200;
			16'h257a: y = 16'h200;
			16'h257b: y = 16'h200;
			16'h257c: y = 16'h200;
			16'h257d: y = 16'h200;
			16'h257e: y = 16'h200;
			16'h257f: y = 16'h200;
			16'h2580: y = 16'h200;
			16'h2581: y = 16'h200;
			16'h2582: y = 16'h200;
			16'h2583: y = 16'h200;
			16'h2584: y = 16'h200;
			16'h2585: y = 16'h200;
			16'h2586: y = 16'h200;
			16'h2587: y = 16'h200;
			16'h2588: y = 16'h200;
			16'h2589: y = 16'h200;
			16'h258a: y = 16'h200;
			16'h258b: y = 16'h200;
			16'h258c: y = 16'h200;
			16'h258d: y = 16'h200;
			16'h258e: y = 16'h200;
			16'h258f: y = 16'h200;
			16'h2590: y = 16'h200;
			16'h2591: y = 16'h200;
			16'h2592: y = 16'h200;
			16'h2593: y = 16'h200;
			16'h2594: y = 16'h200;
			16'h2595: y = 16'h200;
			16'h2596: y = 16'h200;
			16'h2597: y = 16'h200;
			16'h2598: y = 16'h200;
			16'h2599: y = 16'h200;
			16'h259a: y = 16'h200;
			16'h259b: y = 16'h200;
			16'h259c: y = 16'h200;
			16'h259d: y = 16'h200;
			16'h259e: y = 16'h200;
			16'h259f: y = 16'h200;
			16'h25a0: y = 16'h200;
			16'h25a1: y = 16'h200;
			16'h25a2: y = 16'h200;
			16'h25a3: y = 16'h200;
			16'h25a4: y = 16'h200;
			16'h25a5: y = 16'h200;
			16'h25a6: y = 16'h200;
			16'h25a7: y = 16'h200;
			16'h25a8: y = 16'h200;
			16'h25a9: y = 16'h200;
			16'h25aa: y = 16'h200;
			16'h25ab: y = 16'h200;
			16'h25ac: y = 16'h200;
			16'h25ad: y = 16'h200;
			16'h25ae: y = 16'h200;
			16'h25af: y = 16'h200;
			16'h25b0: y = 16'h200;
			16'h25b1: y = 16'h200;
			16'h25b2: y = 16'h200;
			16'h25b3: y = 16'h200;
			16'h25b4: y = 16'h200;
			16'h25b5: y = 16'h200;
			16'h25b6: y = 16'h200;
			16'h25b7: y = 16'h200;
			16'h25b8: y = 16'h200;
			16'h25b9: y = 16'h200;
			16'h25ba: y = 16'h200;
			16'h25bb: y = 16'h200;
			16'h25bc: y = 16'h200;
			16'h25bd: y = 16'h200;
			16'h25be: y = 16'h200;
			16'h25bf: y = 16'h200;
			16'h25c0: y = 16'h200;
			16'h25c1: y = 16'h200;
			16'h25c2: y = 16'h200;
			16'h25c3: y = 16'h200;
			16'h25c4: y = 16'h200;
			16'h25c5: y = 16'h200;
			16'h25c6: y = 16'h200;
			16'h25c7: y = 16'h200;
			16'h25c8: y = 16'h200;
			16'h25c9: y = 16'h200;
			16'h25ca: y = 16'h200;
			16'h25cb: y = 16'h200;
			16'h25cc: y = 16'h200;
			16'h25cd: y = 16'h200;
			16'h25ce: y = 16'h200;
			16'h25cf: y = 16'h200;
			16'h25d0: y = 16'h200;
			16'h25d1: y = 16'h200;
			16'h25d2: y = 16'h200;
			16'h25d3: y = 16'h200;
			16'h25d4: y = 16'h200;
			16'h25d5: y = 16'h200;
			16'h25d6: y = 16'h200;
			16'h25d7: y = 16'h200;
			16'h25d8: y = 16'h200;
			16'h25d9: y = 16'h200;
			16'h25da: y = 16'h200;
			16'h25db: y = 16'h200;
			16'h25dc: y = 16'h200;
			16'h25dd: y = 16'h200;
			16'h25de: y = 16'h200;
			16'h25df: y = 16'h200;
			16'h25e0: y = 16'h200;
			16'h25e1: y = 16'h200;
			16'h25e2: y = 16'h200;
			16'h25e3: y = 16'h200;
			16'h25e4: y = 16'h200;
			16'h25e5: y = 16'h200;
			16'h25e6: y = 16'h200;
			16'h25e7: y = 16'h200;
			16'h25e8: y = 16'h200;
			16'h25e9: y = 16'h200;
			16'h25ea: y = 16'h200;
			16'h25eb: y = 16'h200;
			16'h25ec: y = 16'h200;
			16'h25ed: y = 16'h200;
			16'h25ee: y = 16'h200;
			16'h25ef: y = 16'h200;
			16'h25f0: y = 16'h200;
			16'h25f1: y = 16'h200;
			16'h25f2: y = 16'h200;
			16'h25f3: y = 16'h200;
			16'h25f4: y = 16'h200;
			16'h25f5: y = 16'h200;
			16'h25f6: y = 16'h200;
			16'h25f7: y = 16'h200;
			16'h25f8: y = 16'h200;
			16'h25f9: y = 16'h200;
			16'h25fa: y = 16'h200;
			16'h25fb: y = 16'h200;
			16'h25fc: y = 16'h200;
			16'h25fd: y = 16'h200;
			16'h25fe: y = 16'h200;
			16'h25ff: y = 16'h200;
			16'h2600: y = 16'h200;
			16'h2601: y = 16'h200;
			16'h2602: y = 16'h200;
			16'h2603: y = 16'h200;
			16'h2604: y = 16'h200;
			16'h2605: y = 16'h200;
			16'h2606: y = 16'h200;
			16'h2607: y = 16'h200;
			16'h2608: y = 16'h200;
			16'h2609: y = 16'h200;
			16'h260a: y = 16'h200;
			16'h260b: y = 16'h200;
			16'h260c: y = 16'h200;
			16'h260d: y = 16'h200;
			16'h260e: y = 16'h200;
			16'h260f: y = 16'h200;
			16'h2610: y = 16'h200;
			16'h2611: y = 16'h200;
			16'h2612: y = 16'h200;
			16'h2613: y = 16'h200;
			16'h2614: y = 16'h200;
			16'h2615: y = 16'h200;
			16'h2616: y = 16'h200;
			16'h2617: y = 16'h200;
			16'h2618: y = 16'h200;
			16'h2619: y = 16'h200;
			16'h261a: y = 16'h200;
			16'h261b: y = 16'h200;
			16'h261c: y = 16'h200;
			16'h261d: y = 16'h200;
			16'h261e: y = 16'h200;
			16'h261f: y = 16'h200;
			16'h2620: y = 16'h200;
			16'h2621: y = 16'h200;
			16'h2622: y = 16'h200;
			16'h2623: y = 16'h200;
			16'h2624: y = 16'h200;
			16'h2625: y = 16'h200;
			16'h2626: y = 16'h200;
			16'h2627: y = 16'h200;
			16'h2628: y = 16'h200;
			16'h2629: y = 16'h200;
			16'h262a: y = 16'h200;
			16'h262b: y = 16'h200;
			16'h262c: y = 16'h200;
			16'h262d: y = 16'h200;
			16'h262e: y = 16'h200;
			16'h262f: y = 16'h200;
			16'h2630: y = 16'h200;
			16'h2631: y = 16'h200;
			16'h2632: y = 16'h200;
			16'h2633: y = 16'h200;
			16'h2634: y = 16'h200;
			16'h2635: y = 16'h200;
			16'h2636: y = 16'h200;
			16'h2637: y = 16'h200;
			16'h2638: y = 16'h200;
			16'h2639: y = 16'h200;
			16'h263a: y = 16'h200;
			16'h263b: y = 16'h200;
			16'h263c: y = 16'h200;
			16'h263d: y = 16'h200;
			16'h263e: y = 16'h200;
			16'h263f: y = 16'h200;
			16'h2640: y = 16'h200;
			16'h2641: y = 16'h200;
			16'h2642: y = 16'h200;
			16'h2643: y = 16'h200;
			16'h2644: y = 16'h200;
			16'h2645: y = 16'h200;
			16'h2646: y = 16'h200;
			16'h2647: y = 16'h200;
			16'h2648: y = 16'h200;
			16'h2649: y = 16'h200;
			16'h264a: y = 16'h200;
			16'h264b: y = 16'h200;
			16'h264c: y = 16'h200;
			16'h264d: y = 16'h200;
			16'h264e: y = 16'h200;
			16'h264f: y = 16'h200;
			16'h2650: y = 16'h200;
			16'h2651: y = 16'h200;
			16'h2652: y = 16'h200;
			16'h2653: y = 16'h200;
			16'h2654: y = 16'h200;
			16'h2655: y = 16'h200;
			16'h2656: y = 16'h200;
			16'h2657: y = 16'h200;
			16'h2658: y = 16'h200;
			16'h2659: y = 16'h200;
			16'h265a: y = 16'h200;
			16'h265b: y = 16'h200;
			16'h265c: y = 16'h200;
			16'h265d: y = 16'h200;
			16'h265e: y = 16'h200;
			16'h265f: y = 16'h200;
			16'h2660: y = 16'h200;
			16'h2661: y = 16'h200;
			16'h2662: y = 16'h200;
			16'h2663: y = 16'h200;
			16'h2664: y = 16'h200;
			16'h2665: y = 16'h200;
			16'h2666: y = 16'h200;
			16'h2667: y = 16'h200;
			16'h2668: y = 16'h200;
			16'h2669: y = 16'h200;
			16'h266a: y = 16'h200;
			16'h266b: y = 16'h200;
			16'h266c: y = 16'h200;
			16'h266d: y = 16'h200;
			16'h266e: y = 16'h200;
			16'h266f: y = 16'h200;
			16'h2670: y = 16'h200;
			16'h2671: y = 16'h200;
			16'h2672: y = 16'h200;
			16'h2673: y = 16'h200;
			16'h2674: y = 16'h200;
			16'h2675: y = 16'h200;
			16'h2676: y = 16'h200;
			16'h2677: y = 16'h200;
			16'h2678: y = 16'h200;
			16'h2679: y = 16'h200;
			16'h267a: y = 16'h200;
			16'h267b: y = 16'h200;
			16'h267c: y = 16'h200;
			16'h267d: y = 16'h200;
			16'h267e: y = 16'h200;
			16'h267f: y = 16'h200;
			16'h2680: y = 16'h200;
			16'h2681: y = 16'h200;
			16'h2682: y = 16'h200;
			16'h2683: y = 16'h200;
			16'h2684: y = 16'h200;
			16'h2685: y = 16'h200;
			16'h2686: y = 16'h200;
			16'h2687: y = 16'h200;
			16'h2688: y = 16'h200;
			16'h2689: y = 16'h200;
			16'h268a: y = 16'h200;
			16'h268b: y = 16'h200;
			16'h268c: y = 16'h200;
			16'h268d: y = 16'h200;
			16'h268e: y = 16'h200;
			16'h268f: y = 16'h200;
			16'h2690: y = 16'h200;
			16'h2691: y = 16'h200;
			16'h2692: y = 16'h200;
			16'h2693: y = 16'h200;
			16'h2694: y = 16'h200;
			16'h2695: y = 16'h200;
			16'h2696: y = 16'h200;
			16'h2697: y = 16'h200;
			16'h2698: y = 16'h200;
			16'h2699: y = 16'h200;
			16'h269a: y = 16'h200;
			16'h269b: y = 16'h200;
			16'h269c: y = 16'h200;
			16'h269d: y = 16'h200;
			16'h269e: y = 16'h200;
			16'h269f: y = 16'h200;
			16'h26a0: y = 16'h200;
			16'h26a1: y = 16'h200;
			16'h26a2: y = 16'h200;
			16'h26a3: y = 16'h200;
			16'h26a4: y = 16'h200;
			16'h26a5: y = 16'h200;
			16'h26a6: y = 16'h200;
			16'h26a7: y = 16'h200;
			16'h26a8: y = 16'h200;
			16'h26a9: y = 16'h200;
			16'h26aa: y = 16'h200;
			16'h26ab: y = 16'h200;
			16'h26ac: y = 16'h200;
			16'h26ad: y = 16'h200;
			16'h26ae: y = 16'h200;
			16'h26af: y = 16'h200;
			16'h26b0: y = 16'h200;
			16'h26b1: y = 16'h200;
			16'h26b2: y = 16'h200;
			16'h26b3: y = 16'h200;
			16'h26b4: y = 16'h200;
			16'h26b5: y = 16'h200;
			16'h26b6: y = 16'h200;
			16'h26b7: y = 16'h200;
			16'h26b8: y = 16'h200;
			16'h26b9: y = 16'h200;
			16'h26ba: y = 16'h200;
			16'h26bb: y = 16'h200;
			16'h26bc: y = 16'h200;
			16'h26bd: y = 16'h200;
			16'h26be: y = 16'h200;
			16'h26bf: y = 16'h200;
			16'h26c0: y = 16'h200;
			16'h26c1: y = 16'h200;
			16'h26c2: y = 16'h200;
			16'h26c3: y = 16'h200;
			16'h26c4: y = 16'h200;
			16'h26c5: y = 16'h200;
			16'h26c6: y = 16'h200;
			16'h26c7: y = 16'h200;
			16'h26c8: y = 16'h200;
			16'h26c9: y = 16'h200;
			16'h26ca: y = 16'h200;
			16'h26cb: y = 16'h200;
			16'h26cc: y = 16'h200;
			16'h26cd: y = 16'h200;
			16'h26ce: y = 16'h200;
			16'h26cf: y = 16'h200;
			16'h26d0: y = 16'h200;
			16'h26d1: y = 16'h200;
			16'h26d2: y = 16'h200;
			16'h26d3: y = 16'h200;
			16'h26d4: y = 16'h200;
			16'h26d5: y = 16'h200;
			16'h26d6: y = 16'h200;
			16'h26d7: y = 16'h200;
			16'h26d8: y = 16'h200;
			16'h26d9: y = 16'h200;
			16'h26da: y = 16'h200;
			16'h26db: y = 16'h200;
			16'h26dc: y = 16'h200;
			16'h26dd: y = 16'h200;
			16'h26de: y = 16'h200;
			16'h26df: y = 16'h200;
			16'h26e0: y = 16'h200;
			16'h26e1: y = 16'h200;
			16'h26e2: y = 16'h200;
			16'h26e3: y = 16'h200;
			16'h26e4: y = 16'h200;
			16'h26e5: y = 16'h200;
			16'h26e6: y = 16'h200;
			16'h26e7: y = 16'h200;
			16'h26e8: y = 16'h200;
			16'h26e9: y = 16'h200;
			16'h26ea: y = 16'h200;
			16'h26eb: y = 16'h200;
			16'h26ec: y = 16'h200;
			16'h26ed: y = 16'h200;
			16'h26ee: y = 16'h200;
			16'h26ef: y = 16'h200;
			16'h26f0: y = 16'h200;
			16'h26f1: y = 16'h200;
			16'h26f2: y = 16'h200;
			16'h26f3: y = 16'h200;
			16'h26f4: y = 16'h200;
			16'h26f5: y = 16'h200;
			16'h26f6: y = 16'h200;
			16'h26f7: y = 16'h200;
			16'h26f8: y = 16'h200;
			16'h26f9: y = 16'h200;
			16'h26fa: y = 16'h200;
			16'h26fb: y = 16'h200;
			16'h26fc: y = 16'h200;
			16'h26fd: y = 16'h200;
			16'h26fe: y = 16'h200;
			16'h26ff: y = 16'h200;
			16'h2700: y = 16'h200;
			16'h2701: y = 16'h200;
			16'h2702: y = 16'h200;
			16'h2703: y = 16'h200;
			16'h2704: y = 16'h200;
			16'h2705: y = 16'h200;
			16'h2706: y = 16'h200;
			16'h2707: y = 16'h200;
			16'h2708: y = 16'h200;
			16'h2709: y = 16'h200;
			16'h270a: y = 16'h200;
			16'h270b: y = 16'h200;
			16'h270c: y = 16'h200;
			16'h270d: y = 16'h200;
			16'h270e: y = 16'h200;
			16'h270f: y = 16'h200;
			16'h2710: y = 16'h200;
			16'h2711: y = 16'h200;
			16'h2712: y = 16'h200;
			16'h2713: y = 16'h200;
			16'h2714: y = 16'h200;
			16'h2715: y = 16'h200;
			16'h2716: y = 16'h200;
			16'h2717: y = 16'h200;
			16'h2718: y = 16'h200;
			16'h2719: y = 16'h200;
			16'h271a: y = 16'h200;
			16'h271b: y = 16'h200;
			16'h271c: y = 16'h200;
			16'h271d: y = 16'h200;
			16'h271e: y = 16'h200;
			16'h271f: y = 16'h200;
			16'h2720: y = 16'h200;
			16'h2721: y = 16'h200;
			16'h2722: y = 16'h200;
			16'h2723: y = 16'h200;
			16'h2724: y = 16'h200;
			16'h2725: y = 16'h200;
			16'h2726: y = 16'h200;
			16'h2727: y = 16'h200;
			16'h2728: y = 16'h200;
			16'h2729: y = 16'h200;
			16'h272a: y = 16'h200;
			16'h272b: y = 16'h200;
			16'h272c: y = 16'h200;
			16'h272d: y = 16'h200;
			16'h272e: y = 16'h200;
			16'h272f: y = 16'h200;
			16'h2730: y = 16'h200;
			16'h2731: y = 16'h200;
			16'h2732: y = 16'h200;
			16'h2733: y = 16'h200;
			16'h2734: y = 16'h200;
			16'h2735: y = 16'h200;
			16'h2736: y = 16'h200;
			16'h2737: y = 16'h200;
			16'h2738: y = 16'h200;
			16'h2739: y = 16'h200;
			16'h273a: y = 16'h200;
			16'h273b: y = 16'h200;
			16'h273c: y = 16'h200;
			16'h273d: y = 16'h200;
			16'h273e: y = 16'h200;
			16'h273f: y = 16'h200;
			16'h2740: y = 16'h200;
			16'h2741: y = 16'h200;
			16'h2742: y = 16'h200;
			16'h2743: y = 16'h200;
			16'h2744: y = 16'h200;
			16'h2745: y = 16'h200;
			16'h2746: y = 16'h200;
			16'h2747: y = 16'h200;
			16'h2748: y = 16'h200;
			16'h2749: y = 16'h200;
			16'h274a: y = 16'h200;
			16'h274b: y = 16'h200;
			16'h274c: y = 16'h200;
			16'h274d: y = 16'h200;
			16'h274e: y = 16'h200;
			16'h274f: y = 16'h200;
			16'h2750: y = 16'h200;
			16'h2751: y = 16'h200;
			16'h2752: y = 16'h200;
			16'h2753: y = 16'h200;
			16'h2754: y = 16'h200;
			16'h2755: y = 16'h200;
			16'h2756: y = 16'h200;
			16'h2757: y = 16'h200;
			16'h2758: y = 16'h200;
			16'h2759: y = 16'h200;
			16'h275a: y = 16'h200;
			16'h275b: y = 16'h200;
			16'h275c: y = 16'h200;
			16'h275d: y = 16'h200;
			16'h275e: y = 16'h200;
			16'h275f: y = 16'h200;
			16'h2760: y = 16'h200;
			16'h2761: y = 16'h200;
			16'h2762: y = 16'h200;
			16'h2763: y = 16'h200;
			16'h2764: y = 16'h200;
			16'h2765: y = 16'h200;
			16'h2766: y = 16'h200;
			16'h2767: y = 16'h200;
			16'h2768: y = 16'h200;
			16'h2769: y = 16'h200;
			16'h276a: y = 16'h200;
			16'h276b: y = 16'h200;
			16'h276c: y = 16'h200;
			16'h276d: y = 16'h200;
			16'h276e: y = 16'h200;
			16'h276f: y = 16'h200;
			16'h2770: y = 16'h200;
			16'h2771: y = 16'h200;
			16'h2772: y = 16'h200;
			16'h2773: y = 16'h200;
			16'h2774: y = 16'h200;
			16'h2775: y = 16'h200;
			16'h2776: y = 16'h200;
			16'h2777: y = 16'h200;
			16'h2778: y = 16'h200;
			16'h2779: y = 16'h200;
			16'h277a: y = 16'h200;
			16'h277b: y = 16'h200;
			16'h277c: y = 16'h200;
			16'h277d: y = 16'h200;
			16'h277e: y = 16'h200;
			16'h277f: y = 16'h200;
			16'h2780: y = 16'h200;
			16'h2781: y = 16'h200;
			16'h2782: y = 16'h200;
			16'h2783: y = 16'h200;
			16'h2784: y = 16'h200;
			16'h2785: y = 16'h200;
			16'h2786: y = 16'h200;
			16'h2787: y = 16'h200;
			16'h2788: y = 16'h200;
			16'h2789: y = 16'h200;
			16'h278a: y = 16'h200;
			16'h278b: y = 16'h200;
			16'h278c: y = 16'h200;
			16'h278d: y = 16'h200;
			16'h278e: y = 16'h200;
			16'h278f: y = 16'h200;
			16'h2790: y = 16'h200;
			16'h2791: y = 16'h200;
			16'h2792: y = 16'h200;
			16'h2793: y = 16'h200;
			16'h2794: y = 16'h200;
			16'h2795: y = 16'h200;
			16'h2796: y = 16'h200;
			16'h2797: y = 16'h200;
			16'h2798: y = 16'h200;
			16'h2799: y = 16'h200;
			16'h279a: y = 16'h200;
			16'h279b: y = 16'h200;
			16'h279c: y = 16'h200;
			16'h279d: y = 16'h200;
			16'h279e: y = 16'h200;
			16'h279f: y = 16'h200;
			16'h27a0: y = 16'h200;
			16'h27a1: y = 16'h200;
			16'h27a2: y = 16'h200;
			16'h27a3: y = 16'h200;
			16'h27a4: y = 16'h200;
			16'h27a5: y = 16'h200;
			16'h27a6: y = 16'h200;
			16'h27a7: y = 16'h200;
			16'h27a8: y = 16'h200;
			16'h27a9: y = 16'h200;
			16'h27aa: y = 16'h200;
			16'h27ab: y = 16'h200;
			16'h27ac: y = 16'h200;
			16'h27ad: y = 16'h200;
			16'h27ae: y = 16'h200;
			16'h27af: y = 16'h200;
			16'h27b0: y = 16'h200;
			16'h27b1: y = 16'h200;
			16'h27b2: y = 16'h200;
			16'h27b3: y = 16'h200;
			16'h27b4: y = 16'h200;
			16'h27b5: y = 16'h200;
			16'h27b6: y = 16'h200;
			16'h27b7: y = 16'h200;
			16'h27b8: y = 16'h200;
			16'h27b9: y = 16'h200;
			16'h27ba: y = 16'h200;
			16'h27bb: y = 16'h200;
			16'h27bc: y = 16'h200;
			16'h27bd: y = 16'h200;
			16'h27be: y = 16'h200;
			16'h27bf: y = 16'h200;
			16'h27c0: y = 16'h200;
			16'h27c1: y = 16'h200;
			16'h27c2: y = 16'h200;
			16'h27c3: y = 16'h200;
			16'h27c4: y = 16'h200;
			16'h27c5: y = 16'h200;
			16'h27c6: y = 16'h200;
			16'h27c7: y = 16'h200;
			16'h27c8: y = 16'h200;
			16'h27c9: y = 16'h200;
			16'h27ca: y = 16'h200;
			16'h27cb: y = 16'h200;
			16'h27cc: y = 16'h200;
			16'h27cd: y = 16'h200;
			16'h27ce: y = 16'h200;
			16'h27cf: y = 16'h200;
			16'h27d0: y = 16'h200;
			16'h27d1: y = 16'h200;
			16'h27d2: y = 16'h200;
			16'h27d3: y = 16'h200;
			16'h27d4: y = 16'h200;
			16'h27d5: y = 16'h200;
			16'h27d6: y = 16'h200;
			16'h27d7: y = 16'h200;
			16'h27d8: y = 16'h200;
			16'h27d9: y = 16'h200;
			16'h27da: y = 16'h200;
			16'h27db: y = 16'h200;
			16'h27dc: y = 16'h200;
			16'h27dd: y = 16'h200;
			16'h27de: y = 16'h200;
			16'h27df: y = 16'h200;
			16'h27e0: y = 16'h200;
			16'h27e1: y = 16'h200;
			16'h27e2: y = 16'h200;
			16'h27e3: y = 16'h200;
			16'h27e4: y = 16'h200;
			16'h27e5: y = 16'h200;
			16'h27e6: y = 16'h200;
			16'h27e7: y = 16'h200;
			16'h27e8: y = 16'h200;
			16'h27e9: y = 16'h200;
			16'h27ea: y = 16'h200;
			16'h27eb: y = 16'h200;
			16'h27ec: y = 16'h200;
			16'h27ed: y = 16'h200;
			16'h27ee: y = 16'h200;
			16'h27ef: y = 16'h200;
			16'h27f0: y = 16'h200;
			16'h27f1: y = 16'h200;
			16'h27f2: y = 16'h200;
			16'h27f3: y = 16'h200;
			16'h27f4: y = 16'h200;
			16'h27f5: y = 16'h200;
			16'h27f6: y = 16'h200;
			16'h27f7: y = 16'h200;
			16'h27f8: y = 16'h200;
			16'h27f9: y = 16'h200;
			16'h27fa: y = 16'h200;
			16'h27fb: y = 16'h200;
			16'h27fc: y = 16'h200;
			16'h27fd: y = 16'h200;
			16'h27fe: y = 16'h200;
			16'h27ff: y = 16'h200;
			16'h2800: y = 16'h200;
			16'h2801: y = 16'h200;
			16'h2802: y = 16'h200;
			16'h2803: y = 16'h200;
			16'h2804: y = 16'h200;
			16'h2805: y = 16'h200;
			16'h2806: y = 16'h200;
			16'h2807: y = 16'h200;
			16'h2808: y = 16'h200;
			16'h2809: y = 16'h200;
			16'h280a: y = 16'h200;
			16'h280b: y = 16'h200;
			16'h280c: y = 16'h200;
			16'h280d: y = 16'h200;
			16'h280e: y = 16'h200;
			16'h280f: y = 16'h200;
			16'h2810: y = 16'h200;
			16'h2811: y = 16'h200;
			16'h2812: y = 16'h200;
			16'h2813: y = 16'h200;
			16'h2814: y = 16'h200;
			16'h2815: y = 16'h200;
			16'h2816: y = 16'h200;
			16'h2817: y = 16'h200;
			16'h2818: y = 16'h200;
			16'h2819: y = 16'h200;
			16'h281a: y = 16'h200;
			16'h281b: y = 16'h200;
			16'h281c: y = 16'h200;
			16'h281d: y = 16'h200;
			16'h281e: y = 16'h200;
			16'h281f: y = 16'h200;
			16'h2820: y = 16'h200;
			16'h2821: y = 16'h200;
			16'h2822: y = 16'h200;
			16'h2823: y = 16'h200;
			16'h2824: y = 16'h200;
			16'h2825: y = 16'h200;
			16'h2826: y = 16'h200;
			16'h2827: y = 16'h200;
			16'h2828: y = 16'h200;
			16'h2829: y = 16'h200;
			16'h282a: y = 16'h200;
			16'h282b: y = 16'h200;
			16'h282c: y = 16'h200;
			16'h282d: y = 16'h200;
			16'h282e: y = 16'h200;
			16'h282f: y = 16'h200;
			16'h2830: y = 16'h200;
			16'h2831: y = 16'h200;
			16'h2832: y = 16'h200;
			16'h2833: y = 16'h200;
			16'h2834: y = 16'h200;
			16'h2835: y = 16'h200;
			16'h2836: y = 16'h200;
			16'h2837: y = 16'h200;
			16'h2838: y = 16'h200;
			16'h2839: y = 16'h200;
			16'h283a: y = 16'h200;
			16'h283b: y = 16'h200;
			16'h283c: y = 16'h200;
			16'h283d: y = 16'h200;
			16'h283e: y = 16'h200;
			16'h283f: y = 16'h200;
			16'h2840: y = 16'h200;
			16'h2841: y = 16'h200;
			16'h2842: y = 16'h200;
			16'h2843: y = 16'h200;
			16'h2844: y = 16'h200;
			16'h2845: y = 16'h200;
			16'h2846: y = 16'h200;
			16'h2847: y = 16'h200;
			16'h2848: y = 16'h200;
			16'h2849: y = 16'h200;
			16'h284a: y = 16'h200;
			16'h284b: y = 16'h200;
			16'h284c: y = 16'h200;
			16'h284d: y = 16'h200;
			16'h284e: y = 16'h200;
			16'h284f: y = 16'h200;
			16'h2850: y = 16'h200;
			16'h2851: y = 16'h200;
			16'h2852: y = 16'h200;
			16'h2853: y = 16'h200;
			16'h2854: y = 16'h200;
			16'h2855: y = 16'h200;
			16'h2856: y = 16'h200;
			16'h2857: y = 16'h200;
			16'h2858: y = 16'h200;
			16'h2859: y = 16'h200;
			16'h285a: y = 16'h200;
			16'h285b: y = 16'h200;
			16'h285c: y = 16'h200;
			16'h285d: y = 16'h200;
			16'h285e: y = 16'h200;
			16'h285f: y = 16'h200;
			16'h2860: y = 16'h200;
			16'h2861: y = 16'h200;
			16'h2862: y = 16'h200;
			16'h2863: y = 16'h200;
			16'h2864: y = 16'h200;
			16'h2865: y = 16'h200;
			16'h2866: y = 16'h200;
			16'h2867: y = 16'h200;
			16'h2868: y = 16'h200;
			16'h2869: y = 16'h200;
			16'h286a: y = 16'h200;
			16'h286b: y = 16'h200;
			16'h286c: y = 16'h200;
			16'h286d: y = 16'h200;
			16'h286e: y = 16'h200;
			16'h286f: y = 16'h200;
			16'h2870: y = 16'h200;
			16'h2871: y = 16'h200;
			16'h2872: y = 16'h200;
			16'h2873: y = 16'h200;
			16'h2874: y = 16'h200;
			16'h2875: y = 16'h200;
			16'h2876: y = 16'h200;
			16'h2877: y = 16'h200;
			16'h2878: y = 16'h200;
			16'h2879: y = 16'h200;
			16'h287a: y = 16'h200;
			16'h287b: y = 16'h200;
			16'h287c: y = 16'h200;
			16'h287d: y = 16'h200;
			16'h287e: y = 16'h200;
			16'h287f: y = 16'h200;
			16'h2880: y = 16'h200;
			16'h2881: y = 16'h200;
			16'h2882: y = 16'h200;
			16'h2883: y = 16'h200;
			16'h2884: y = 16'h200;
			16'h2885: y = 16'h200;
			16'h2886: y = 16'h200;
			16'h2887: y = 16'h200;
			16'h2888: y = 16'h200;
			16'h2889: y = 16'h200;
			16'h288a: y = 16'h200;
			16'h288b: y = 16'h200;
			16'h288c: y = 16'h200;
			16'h288d: y = 16'h200;
			16'h288e: y = 16'h200;
			16'h288f: y = 16'h200;
			16'h2890: y = 16'h200;
			16'h2891: y = 16'h200;
			16'h2892: y = 16'h200;
			16'h2893: y = 16'h200;
			16'h2894: y = 16'h200;
			16'h2895: y = 16'h200;
			16'h2896: y = 16'h200;
			16'h2897: y = 16'h200;
			16'h2898: y = 16'h200;
			16'h2899: y = 16'h200;
			16'h289a: y = 16'h200;
			16'h289b: y = 16'h200;
			16'h289c: y = 16'h200;
			16'h289d: y = 16'h200;
			16'h289e: y = 16'h200;
			16'h289f: y = 16'h200;
			16'h28a0: y = 16'h200;
			16'h28a1: y = 16'h200;
			16'h28a2: y = 16'h200;
			16'h28a3: y = 16'h200;
			16'h28a4: y = 16'h200;
			16'h28a5: y = 16'h200;
			16'h28a6: y = 16'h200;
			16'h28a7: y = 16'h200;
			16'h28a8: y = 16'h200;
			16'h28a9: y = 16'h200;
			16'h28aa: y = 16'h200;
			16'h28ab: y = 16'h200;
			16'h28ac: y = 16'h200;
			16'h28ad: y = 16'h200;
			16'h28ae: y = 16'h200;
			16'h28af: y = 16'h200;
			16'h28b0: y = 16'h200;
			16'h28b1: y = 16'h200;
			16'h28b2: y = 16'h200;
			16'h28b3: y = 16'h200;
			16'h28b4: y = 16'h200;
			16'h28b5: y = 16'h200;
			16'h28b6: y = 16'h200;
			16'h28b7: y = 16'h200;
			16'h28b8: y = 16'h200;
			16'h28b9: y = 16'h200;
			16'h28ba: y = 16'h200;
			16'h28bb: y = 16'h200;
			16'h28bc: y = 16'h200;
			16'h28bd: y = 16'h200;
			16'h28be: y = 16'h200;
			16'h28bf: y = 16'h200;
			16'h28c0: y = 16'h200;
			16'h28c1: y = 16'h200;
			16'h28c2: y = 16'h200;
			16'h28c3: y = 16'h200;
			16'h28c4: y = 16'h200;
			16'h28c5: y = 16'h200;
			16'h28c6: y = 16'h200;
			16'h28c7: y = 16'h200;
			16'h28c8: y = 16'h200;
			16'h28c9: y = 16'h200;
			16'h28ca: y = 16'h200;
			16'h28cb: y = 16'h200;
			16'h28cc: y = 16'h200;
			16'h28cd: y = 16'h200;
			16'h28ce: y = 16'h200;
			16'h28cf: y = 16'h200;
			16'h28d0: y = 16'h200;
			16'h28d1: y = 16'h200;
			16'h28d2: y = 16'h200;
			16'h28d3: y = 16'h200;
			16'h28d4: y = 16'h200;
			16'h28d5: y = 16'h200;
			16'h28d6: y = 16'h200;
			16'h28d7: y = 16'h200;
			16'h28d8: y = 16'h200;
			16'h28d9: y = 16'h200;
			16'h28da: y = 16'h200;
			16'h28db: y = 16'h200;
			16'h28dc: y = 16'h200;
			16'h28dd: y = 16'h200;
			16'h28de: y = 16'h200;
			16'h28df: y = 16'h200;
			16'h28e0: y = 16'h200;
			16'h28e1: y = 16'h200;
			16'h28e2: y = 16'h200;
			16'h28e3: y = 16'h200;
			16'h28e4: y = 16'h200;
			16'h28e5: y = 16'h200;
			16'h28e6: y = 16'h200;
			16'h28e7: y = 16'h200;
			16'h28e8: y = 16'h200;
			16'h28e9: y = 16'h200;
			16'h28ea: y = 16'h200;
			16'h28eb: y = 16'h200;
			16'h28ec: y = 16'h200;
			16'h28ed: y = 16'h200;
			16'h28ee: y = 16'h200;
			16'h28ef: y = 16'h200;
			16'h28f0: y = 16'h200;
			16'h28f1: y = 16'h200;
			16'h28f2: y = 16'h200;
			16'h28f3: y = 16'h200;
			16'h28f4: y = 16'h200;
			16'h28f5: y = 16'h200;
			16'h28f6: y = 16'h200;
			16'h28f7: y = 16'h200;
			16'h28f8: y = 16'h200;
			16'h28f9: y = 16'h200;
			16'h28fa: y = 16'h200;
			16'h28fb: y = 16'h200;
			16'h28fc: y = 16'h200;
			16'h28fd: y = 16'h200;
			16'h28fe: y = 16'h200;
			16'h28ff: y = 16'h200;
			16'h2900: y = 16'h200;
			16'h2901: y = 16'h200;
			16'h2902: y = 16'h200;
			16'h2903: y = 16'h200;
			16'h2904: y = 16'h200;
			16'h2905: y = 16'h200;
			16'h2906: y = 16'h200;
			16'h2907: y = 16'h200;
			16'h2908: y = 16'h200;
			16'h2909: y = 16'h200;
			16'h290a: y = 16'h200;
			16'h290b: y = 16'h200;
			16'h290c: y = 16'h200;
			16'h290d: y = 16'h200;
			16'h290e: y = 16'h200;
			16'h290f: y = 16'h200;
			16'h2910: y = 16'h200;
			16'h2911: y = 16'h200;
			16'h2912: y = 16'h200;
			16'h2913: y = 16'h200;
			16'h2914: y = 16'h200;
			16'h2915: y = 16'h200;
			16'h2916: y = 16'h200;
			16'h2917: y = 16'h200;
			16'h2918: y = 16'h200;
			16'h2919: y = 16'h200;
			16'h291a: y = 16'h200;
			16'h291b: y = 16'h200;
			16'h291c: y = 16'h200;
			16'h291d: y = 16'h200;
			16'h291e: y = 16'h200;
			16'h291f: y = 16'h200;
			16'h2920: y = 16'h200;
			16'h2921: y = 16'h200;
			16'h2922: y = 16'h200;
			16'h2923: y = 16'h200;
			16'h2924: y = 16'h200;
			16'h2925: y = 16'h200;
			16'h2926: y = 16'h200;
			16'h2927: y = 16'h200;
			16'h2928: y = 16'h200;
			16'h2929: y = 16'h200;
			16'h292a: y = 16'h200;
			16'h292b: y = 16'h200;
			16'h292c: y = 16'h200;
			16'h292d: y = 16'h200;
			16'h292e: y = 16'h200;
			16'h292f: y = 16'h200;
			16'h2930: y = 16'h200;
			16'h2931: y = 16'h200;
			16'h2932: y = 16'h200;
			16'h2933: y = 16'h200;
			16'h2934: y = 16'h200;
			16'h2935: y = 16'h200;
			16'h2936: y = 16'h200;
			16'h2937: y = 16'h200;
			16'h2938: y = 16'h200;
			16'h2939: y = 16'h200;
			16'h293a: y = 16'h200;
			16'h293b: y = 16'h200;
			16'h293c: y = 16'h200;
			16'h293d: y = 16'h200;
			16'h293e: y = 16'h200;
			16'h293f: y = 16'h200;
			16'h2940: y = 16'h200;
			16'h2941: y = 16'h200;
			16'h2942: y = 16'h200;
			16'h2943: y = 16'h200;
			16'h2944: y = 16'h200;
			16'h2945: y = 16'h200;
			16'h2946: y = 16'h200;
			16'h2947: y = 16'h200;
			16'h2948: y = 16'h200;
			16'h2949: y = 16'h200;
			16'h294a: y = 16'h200;
			16'h294b: y = 16'h200;
			16'h294c: y = 16'h200;
			16'h294d: y = 16'h200;
			16'h294e: y = 16'h200;
			16'h294f: y = 16'h200;
			16'h2950: y = 16'h200;
			16'h2951: y = 16'h200;
			16'h2952: y = 16'h200;
			16'h2953: y = 16'h200;
			16'h2954: y = 16'h200;
			16'h2955: y = 16'h200;
			16'h2956: y = 16'h200;
			16'h2957: y = 16'h200;
			16'h2958: y = 16'h200;
			16'h2959: y = 16'h200;
			16'h295a: y = 16'h200;
			16'h295b: y = 16'h200;
			16'h295c: y = 16'h200;
			16'h295d: y = 16'h200;
			16'h295e: y = 16'h200;
			16'h295f: y = 16'h200;
			16'h2960: y = 16'h200;
			16'h2961: y = 16'h200;
			16'h2962: y = 16'h200;
			16'h2963: y = 16'h200;
			16'h2964: y = 16'h200;
			16'h2965: y = 16'h200;
			16'h2966: y = 16'h200;
			16'h2967: y = 16'h200;
			16'h2968: y = 16'h200;
			16'h2969: y = 16'h200;
			16'h296a: y = 16'h200;
			16'h296b: y = 16'h200;
			16'h296c: y = 16'h200;
			16'h296d: y = 16'h200;
			16'h296e: y = 16'h200;
			16'h296f: y = 16'h200;
			16'h2970: y = 16'h200;
			16'h2971: y = 16'h200;
			16'h2972: y = 16'h200;
			16'h2973: y = 16'h200;
			16'h2974: y = 16'h200;
			16'h2975: y = 16'h200;
			16'h2976: y = 16'h200;
			16'h2977: y = 16'h200;
			16'h2978: y = 16'h200;
			16'h2979: y = 16'h200;
			16'h297a: y = 16'h200;
			16'h297b: y = 16'h200;
			16'h297c: y = 16'h200;
			16'h297d: y = 16'h200;
			16'h297e: y = 16'h200;
			16'h297f: y = 16'h200;
			16'h2980: y = 16'h200;
			16'h2981: y = 16'h200;
			16'h2982: y = 16'h200;
			16'h2983: y = 16'h200;
			16'h2984: y = 16'h200;
			16'h2985: y = 16'h200;
			16'h2986: y = 16'h200;
			16'h2987: y = 16'h200;
			16'h2988: y = 16'h200;
			16'h2989: y = 16'h200;
			16'h298a: y = 16'h200;
			16'h298b: y = 16'h200;
			16'h298c: y = 16'h200;
			16'h298d: y = 16'h200;
			16'h298e: y = 16'h200;
			16'h298f: y = 16'h200;
			16'h2990: y = 16'h200;
			16'h2991: y = 16'h200;
			16'h2992: y = 16'h200;
			16'h2993: y = 16'h200;
			16'h2994: y = 16'h200;
			16'h2995: y = 16'h200;
			16'h2996: y = 16'h200;
			16'h2997: y = 16'h200;
			16'h2998: y = 16'h200;
			16'h2999: y = 16'h200;
			16'h299a: y = 16'h200;
			16'h299b: y = 16'h200;
			16'h299c: y = 16'h200;
			16'h299d: y = 16'h200;
			16'h299e: y = 16'h200;
			16'h299f: y = 16'h200;
			16'h29a0: y = 16'h200;
			16'h29a1: y = 16'h200;
			16'h29a2: y = 16'h200;
			16'h29a3: y = 16'h200;
			16'h29a4: y = 16'h200;
			16'h29a5: y = 16'h200;
			16'h29a6: y = 16'h200;
			16'h29a7: y = 16'h200;
			16'h29a8: y = 16'h200;
			16'h29a9: y = 16'h200;
			16'h29aa: y = 16'h200;
			16'h29ab: y = 16'h200;
			16'h29ac: y = 16'h200;
			16'h29ad: y = 16'h200;
			16'h29ae: y = 16'h200;
			16'h29af: y = 16'h200;
			16'h29b0: y = 16'h200;
			16'h29b1: y = 16'h200;
			16'h29b2: y = 16'h200;
			16'h29b3: y = 16'h200;
			16'h29b4: y = 16'h200;
			16'h29b5: y = 16'h200;
			16'h29b6: y = 16'h200;
			16'h29b7: y = 16'h200;
			16'h29b8: y = 16'h200;
			16'h29b9: y = 16'h200;
			16'h29ba: y = 16'h200;
			16'h29bb: y = 16'h200;
			16'h29bc: y = 16'h200;
			16'h29bd: y = 16'h200;
			16'h29be: y = 16'h200;
			16'h29bf: y = 16'h200;
			16'h29c0: y = 16'h200;
			16'h29c1: y = 16'h200;
			16'h29c2: y = 16'h200;
			16'h29c3: y = 16'h200;
			16'h29c4: y = 16'h200;
			16'h29c5: y = 16'h200;
			16'h29c6: y = 16'h200;
			16'h29c7: y = 16'h200;
			16'h29c8: y = 16'h200;
			16'h29c9: y = 16'h200;
			16'h29ca: y = 16'h200;
			16'h29cb: y = 16'h200;
			16'h29cc: y = 16'h200;
			16'h29cd: y = 16'h200;
			16'h29ce: y = 16'h200;
			16'h29cf: y = 16'h200;
			16'h29d0: y = 16'h200;
			16'h29d1: y = 16'h200;
			16'h29d2: y = 16'h200;
			16'h29d3: y = 16'h200;
			16'h29d4: y = 16'h200;
			16'h29d5: y = 16'h200;
			16'h29d6: y = 16'h200;
			16'h29d7: y = 16'h200;
			16'h29d8: y = 16'h200;
			16'h29d9: y = 16'h200;
			16'h29da: y = 16'h200;
			16'h29db: y = 16'h200;
			16'h29dc: y = 16'h200;
			16'h29dd: y = 16'h200;
			16'h29de: y = 16'h200;
			16'h29df: y = 16'h200;
			16'h29e0: y = 16'h200;
			16'h29e1: y = 16'h200;
			16'h29e2: y = 16'h200;
			16'h29e3: y = 16'h200;
			16'h29e4: y = 16'h200;
			16'h29e5: y = 16'h200;
			16'h29e6: y = 16'h200;
			16'h29e7: y = 16'h200;
			16'h29e8: y = 16'h200;
			16'h29e9: y = 16'h200;
			16'h29ea: y = 16'h200;
			16'h29eb: y = 16'h200;
			16'h29ec: y = 16'h200;
			16'h29ed: y = 16'h200;
			16'h29ee: y = 16'h200;
			16'h29ef: y = 16'h200;
			16'h29f0: y = 16'h200;
			16'h29f1: y = 16'h200;
			16'h29f2: y = 16'h200;
			16'h29f3: y = 16'h200;
			16'h29f4: y = 16'h200;
			16'h29f5: y = 16'h200;
			16'h29f6: y = 16'h200;
			16'h29f7: y = 16'h200;
			16'h29f8: y = 16'h200;
			16'h29f9: y = 16'h200;
			16'h29fa: y = 16'h200;
			16'h29fb: y = 16'h200;
			16'h29fc: y = 16'h200;
			16'h29fd: y = 16'h200;
			16'h29fe: y = 16'h200;
			16'h29ff: y = 16'h200;
			16'h2a00: y = 16'h200;
			16'h2a01: y = 16'h200;
			16'h2a02: y = 16'h200;
			16'h2a03: y = 16'h200;
			16'h2a04: y = 16'h200;
			16'h2a05: y = 16'h200;
			16'h2a06: y = 16'h200;
			16'h2a07: y = 16'h200;
			16'h2a08: y = 16'h200;
			16'h2a09: y = 16'h200;
			16'h2a0a: y = 16'h200;
			16'h2a0b: y = 16'h200;
			16'h2a0c: y = 16'h200;
			16'h2a0d: y = 16'h200;
			16'h2a0e: y = 16'h200;
			16'h2a0f: y = 16'h200;
			16'h2a10: y = 16'h200;
			16'h2a11: y = 16'h200;
			16'h2a12: y = 16'h200;
			16'h2a13: y = 16'h200;
			16'h2a14: y = 16'h200;
			16'h2a15: y = 16'h200;
			16'h2a16: y = 16'h200;
			16'h2a17: y = 16'h200;
			16'h2a18: y = 16'h200;
			16'h2a19: y = 16'h200;
			16'h2a1a: y = 16'h200;
			16'h2a1b: y = 16'h200;
			16'h2a1c: y = 16'h200;
			16'h2a1d: y = 16'h200;
			16'h2a1e: y = 16'h200;
			16'h2a1f: y = 16'h200;
			16'h2a20: y = 16'h200;
			16'h2a21: y = 16'h200;
			16'h2a22: y = 16'h200;
			16'h2a23: y = 16'h200;
			16'h2a24: y = 16'h200;
			16'h2a25: y = 16'h200;
			16'h2a26: y = 16'h200;
			16'h2a27: y = 16'h200;
			16'h2a28: y = 16'h200;
			16'h2a29: y = 16'h200;
			16'h2a2a: y = 16'h200;
			16'h2a2b: y = 16'h200;
			16'h2a2c: y = 16'h200;
			16'h2a2d: y = 16'h200;
			16'h2a2e: y = 16'h200;
			16'h2a2f: y = 16'h200;
			16'h2a30: y = 16'h200;
			16'h2a31: y = 16'h200;
			16'h2a32: y = 16'h200;
			16'h2a33: y = 16'h200;
			16'h2a34: y = 16'h200;
			16'h2a35: y = 16'h200;
			16'h2a36: y = 16'h200;
			16'h2a37: y = 16'h200;
			16'h2a38: y = 16'h200;
			16'h2a39: y = 16'h200;
			16'h2a3a: y = 16'h200;
			16'h2a3b: y = 16'h200;
			16'h2a3c: y = 16'h200;
			16'h2a3d: y = 16'h200;
			16'h2a3e: y = 16'h200;
			16'h2a3f: y = 16'h200;
			16'h2a40: y = 16'h200;
			16'h2a41: y = 16'h200;
			16'h2a42: y = 16'h200;
			16'h2a43: y = 16'h200;
			16'h2a44: y = 16'h200;
			16'h2a45: y = 16'h200;
			16'h2a46: y = 16'h200;
			16'h2a47: y = 16'h200;
			16'h2a48: y = 16'h200;
			16'h2a49: y = 16'h200;
			16'h2a4a: y = 16'h200;
			16'h2a4b: y = 16'h200;
			16'h2a4c: y = 16'h200;
			16'h2a4d: y = 16'h200;
			16'h2a4e: y = 16'h200;
			16'h2a4f: y = 16'h200;
			16'h2a50: y = 16'h200;
			16'h2a51: y = 16'h200;
			16'h2a52: y = 16'h200;
			16'h2a53: y = 16'h200;
			16'h2a54: y = 16'h200;
			16'h2a55: y = 16'h200;
			16'h2a56: y = 16'h200;
			16'h2a57: y = 16'h200;
			16'h2a58: y = 16'h200;
			16'h2a59: y = 16'h200;
			16'h2a5a: y = 16'h200;
			16'h2a5b: y = 16'h200;
			16'h2a5c: y = 16'h200;
			16'h2a5d: y = 16'h200;
			16'h2a5e: y = 16'h200;
			16'h2a5f: y = 16'h200;
			16'h2a60: y = 16'h200;
			16'h2a61: y = 16'h200;
			16'h2a62: y = 16'h200;
			16'h2a63: y = 16'h200;
			16'h2a64: y = 16'h200;
			16'h2a65: y = 16'h200;
			16'h2a66: y = 16'h200;
			16'h2a67: y = 16'h200;
			16'h2a68: y = 16'h200;
			16'h2a69: y = 16'h200;
			16'h2a6a: y = 16'h200;
			16'h2a6b: y = 16'h200;
			16'h2a6c: y = 16'h200;
			16'h2a6d: y = 16'h200;
			16'h2a6e: y = 16'h200;
			16'h2a6f: y = 16'h200;
			16'h2a70: y = 16'h200;
			16'h2a71: y = 16'h200;
			16'h2a72: y = 16'h200;
			16'h2a73: y = 16'h200;
			16'h2a74: y = 16'h200;
			16'h2a75: y = 16'h200;
			16'h2a76: y = 16'h200;
			16'h2a77: y = 16'h200;
			16'h2a78: y = 16'h200;
			16'h2a79: y = 16'h200;
			16'h2a7a: y = 16'h200;
			16'h2a7b: y = 16'h200;
			16'h2a7c: y = 16'h200;
			16'h2a7d: y = 16'h200;
			16'h2a7e: y = 16'h200;
			16'h2a7f: y = 16'h200;
			16'h2a80: y = 16'h200;
			16'h2a81: y = 16'h200;
			16'h2a82: y = 16'h200;
			16'h2a83: y = 16'h200;
			16'h2a84: y = 16'h200;
			16'h2a85: y = 16'h200;
			16'h2a86: y = 16'h200;
			16'h2a87: y = 16'h200;
			16'h2a88: y = 16'h200;
			16'h2a89: y = 16'h200;
			16'h2a8a: y = 16'h200;
			16'h2a8b: y = 16'h200;
			16'h2a8c: y = 16'h200;
			16'h2a8d: y = 16'h200;
			16'h2a8e: y = 16'h200;
			16'h2a8f: y = 16'h200;
			16'h2a90: y = 16'h200;
			16'h2a91: y = 16'h200;
			16'h2a92: y = 16'h200;
			16'h2a93: y = 16'h200;
			16'h2a94: y = 16'h200;
			16'h2a95: y = 16'h200;
			16'h2a96: y = 16'h200;
			16'h2a97: y = 16'h200;
			16'h2a98: y = 16'h200;
			16'h2a99: y = 16'h200;
			16'h2a9a: y = 16'h200;
			16'h2a9b: y = 16'h200;
			16'h2a9c: y = 16'h200;
			16'h2a9d: y = 16'h200;
			16'h2a9e: y = 16'h200;
			16'h2a9f: y = 16'h200;
			16'h2aa0: y = 16'h200;
			16'h2aa1: y = 16'h200;
			16'h2aa2: y = 16'h200;
			16'h2aa3: y = 16'h200;
			16'h2aa4: y = 16'h200;
			16'h2aa5: y = 16'h200;
			16'h2aa6: y = 16'h200;
			16'h2aa7: y = 16'h200;
			16'h2aa8: y = 16'h200;
			16'h2aa9: y = 16'h200;
			16'h2aaa: y = 16'h200;
			16'h2aab: y = 16'h200;
			16'h2aac: y = 16'h200;
			16'h2aad: y = 16'h200;
			16'h2aae: y = 16'h200;
			16'h2aaf: y = 16'h200;
			16'h2ab0: y = 16'h200;
			16'h2ab1: y = 16'h200;
			16'h2ab2: y = 16'h200;
			16'h2ab3: y = 16'h200;
			16'h2ab4: y = 16'h200;
			16'h2ab5: y = 16'h200;
			16'h2ab6: y = 16'h200;
			16'h2ab7: y = 16'h200;
			16'h2ab8: y = 16'h200;
			16'h2ab9: y = 16'h200;
			16'h2aba: y = 16'h200;
			16'h2abb: y = 16'h200;
			16'h2abc: y = 16'h200;
			16'h2abd: y = 16'h200;
			16'h2abe: y = 16'h200;
			16'h2abf: y = 16'h200;
			16'h2ac0: y = 16'h200;
			16'h2ac1: y = 16'h200;
			16'h2ac2: y = 16'h200;
			16'h2ac3: y = 16'h200;
			16'h2ac4: y = 16'h200;
			16'h2ac5: y = 16'h200;
			16'h2ac6: y = 16'h200;
			16'h2ac7: y = 16'h200;
			16'h2ac8: y = 16'h200;
			16'h2ac9: y = 16'h200;
			16'h2aca: y = 16'h200;
			16'h2acb: y = 16'h200;
			16'h2acc: y = 16'h200;
			16'h2acd: y = 16'h200;
			16'h2ace: y = 16'h200;
			16'h2acf: y = 16'h200;
			16'h2ad0: y = 16'h200;
			16'h2ad1: y = 16'h200;
			16'h2ad2: y = 16'h200;
			16'h2ad3: y = 16'h200;
			16'h2ad4: y = 16'h200;
			16'h2ad5: y = 16'h200;
			16'h2ad6: y = 16'h200;
			16'h2ad7: y = 16'h200;
			16'h2ad8: y = 16'h200;
			16'h2ad9: y = 16'h200;
			16'h2ada: y = 16'h200;
			16'h2adb: y = 16'h200;
			16'h2adc: y = 16'h200;
			16'h2add: y = 16'h200;
			16'h2ade: y = 16'h200;
			16'h2adf: y = 16'h200;
			16'h2ae0: y = 16'h200;
			16'h2ae1: y = 16'h200;
			16'h2ae2: y = 16'h200;
			16'h2ae3: y = 16'h200;
			16'h2ae4: y = 16'h200;
			16'h2ae5: y = 16'h200;
			16'h2ae6: y = 16'h200;
			16'h2ae7: y = 16'h200;
			16'h2ae8: y = 16'h200;
			16'h2ae9: y = 16'h200;
			16'h2aea: y = 16'h200;
			16'h2aeb: y = 16'h200;
			16'h2aec: y = 16'h200;
			16'h2aed: y = 16'h200;
			16'h2aee: y = 16'h200;
			16'h2aef: y = 16'h200;
			16'h2af0: y = 16'h200;
			16'h2af1: y = 16'h200;
			16'h2af2: y = 16'h200;
			16'h2af3: y = 16'h200;
			16'h2af4: y = 16'h200;
			16'h2af5: y = 16'h200;
			16'h2af6: y = 16'h200;
			16'h2af7: y = 16'h200;
			16'h2af8: y = 16'h200;
			16'h2af9: y = 16'h200;
			16'h2afa: y = 16'h200;
			16'h2afb: y = 16'h200;
			16'h2afc: y = 16'h200;
			16'h2afd: y = 16'h200;
			16'h2afe: y = 16'h200;
			16'h2aff: y = 16'h200;
			16'h2b00: y = 16'h200;
			16'h2b01: y = 16'h200;
			16'h2b02: y = 16'h200;
			16'h2b03: y = 16'h200;
			16'h2b04: y = 16'h200;
			16'h2b05: y = 16'h200;
			16'h2b06: y = 16'h200;
			16'h2b07: y = 16'h200;
			16'h2b08: y = 16'h200;
			16'h2b09: y = 16'h200;
			16'h2b0a: y = 16'h200;
			16'h2b0b: y = 16'h200;
			16'h2b0c: y = 16'h200;
			16'h2b0d: y = 16'h200;
			16'h2b0e: y = 16'h200;
			16'h2b0f: y = 16'h200;
			16'h2b10: y = 16'h200;
			16'h2b11: y = 16'h200;
			16'h2b12: y = 16'h200;
			16'h2b13: y = 16'h200;
			16'h2b14: y = 16'h200;
			16'h2b15: y = 16'h200;
			16'h2b16: y = 16'h200;
			16'h2b17: y = 16'h200;
			16'h2b18: y = 16'h200;
			16'h2b19: y = 16'h200;
			16'h2b1a: y = 16'h200;
			16'h2b1b: y = 16'h200;
			16'h2b1c: y = 16'h200;
			16'h2b1d: y = 16'h200;
			16'h2b1e: y = 16'h200;
			16'h2b1f: y = 16'h200;
			16'h2b20: y = 16'h200;
			16'h2b21: y = 16'h200;
			16'h2b22: y = 16'h200;
			16'h2b23: y = 16'h200;
			16'h2b24: y = 16'h200;
			16'h2b25: y = 16'h200;
			16'h2b26: y = 16'h200;
			16'h2b27: y = 16'h200;
			16'h2b28: y = 16'h200;
			16'h2b29: y = 16'h200;
			16'h2b2a: y = 16'h200;
			16'h2b2b: y = 16'h200;
			16'h2b2c: y = 16'h200;
			16'h2b2d: y = 16'h200;
			16'h2b2e: y = 16'h200;
			16'h2b2f: y = 16'h200;
			16'h2b30: y = 16'h200;
			16'h2b31: y = 16'h200;
			16'h2b32: y = 16'h200;
			16'h2b33: y = 16'h200;
			16'h2b34: y = 16'h200;
			16'h2b35: y = 16'h200;
			16'h2b36: y = 16'h200;
			16'h2b37: y = 16'h200;
			16'h2b38: y = 16'h200;
			16'h2b39: y = 16'h200;
			16'h2b3a: y = 16'h200;
			16'h2b3b: y = 16'h200;
			16'h2b3c: y = 16'h200;
			16'h2b3d: y = 16'h200;
			16'h2b3e: y = 16'h200;
			16'h2b3f: y = 16'h200;
			16'h2b40: y = 16'h200;
			16'h2b41: y = 16'h200;
			16'h2b42: y = 16'h200;
			16'h2b43: y = 16'h200;
			16'h2b44: y = 16'h200;
			16'h2b45: y = 16'h200;
			16'h2b46: y = 16'h200;
			16'h2b47: y = 16'h200;
			16'h2b48: y = 16'h200;
			16'h2b49: y = 16'h200;
			16'h2b4a: y = 16'h200;
			16'h2b4b: y = 16'h200;
			16'h2b4c: y = 16'h200;
			16'h2b4d: y = 16'h200;
			16'h2b4e: y = 16'h200;
			16'h2b4f: y = 16'h200;
			16'h2b50: y = 16'h200;
			16'h2b51: y = 16'h200;
			16'h2b52: y = 16'h200;
			16'h2b53: y = 16'h200;
			16'h2b54: y = 16'h200;
			16'h2b55: y = 16'h200;
			16'h2b56: y = 16'h200;
			16'h2b57: y = 16'h200;
			16'h2b58: y = 16'h200;
			16'h2b59: y = 16'h200;
			16'h2b5a: y = 16'h200;
			16'h2b5b: y = 16'h200;
			16'h2b5c: y = 16'h200;
			16'h2b5d: y = 16'h200;
			16'h2b5e: y = 16'h200;
			16'h2b5f: y = 16'h200;
			16'h2b60: y = 16'h200;
			16'h2b61: y = 16'h200;
			16'h2b62: y = 16'h200;
			16'h2b63: y = 16'h200;
			16'h2b64: y = 16'h200;
			16'h2b65: y = 16'h200;
			16'h2b66: y = 16'h200;
			16'h2b67: y = 16'h200;
			16'h2b68: y = 16'h200;
			16'h2b69: y = 16'h200;
			16'h2b6a: y = 16'h200;
			16'h2b6b: y = 16'h200;
			16'h2b6c: y = 16'h200;
			16'h2b6d: y = 16'h200;
			16'h2b6e: y = 16'h200;
			16'h2b6f: y = 16'h200;
			16'h2b70: y = 16'h200;
			16'h2b71: y = 16'h200;
			16'h2b72: y = 16'h200;
			16'h2b73: y = 16'h200;
			16'h2b74: y = 16'h200;
			16'h2b75: y = 16'h200;
			16'h2b76: y = 16'h200;
			16'h2b77: y = 16'h200;
			16'h2b78: y = 16'h200;
			16'h2b79: y = 16'h200;
			16'h2b7a: y = 16'h200;
			16'h2b7b: y = 16'h200;
			16'h2b7c: y = 16'h200;
			16'h2b7d: y = 16'h200;
			16'h2b7e: y = 16'h200;
			16'h2b7f: y = 16'h200;
			16'h2b80: y = 16'h200;
			16'h2b81: y = 16'h200;
			16'h2b82: y = 16'h200;
			16'h2b83: y = 16'h200;
			16'h2b84: y = 16'h200;
			16'h2b85: y = 16'h200;
			16'h2b86: y = 16'h200;
			16'h2b87: y = 16'h200;
			16'h2b88: y = 16'h200;
			16'h2b89: y = 16'h200;
			16'h2b8a: y = 16'h200;
			16'h2b8b: y = 16'h200;
			16'h2b8c: y = 16'h200;
			16'h2b8d: y = 16'h200;
			16'h2b8e: y = 16'h200;
			16'h2b8f: y = 16'h200;
			16'h2b90: y = 16'h200;
			16'h2b91: y = 16'h200;
			16'h2b92: y = 16'h200;
			16'h2b93: y = 16'h200;
			16'h2b94: y = 16'h200;
			16'h2b95: y = 16'h200;
			16'h2b96: y = 16'h200;
			16'h2b97: y = 16'h200;
			16'h2b98: y = 16'h200;
			16'h2b99: y = 16'h200;
			16'h2b9a: y = 16'h200;
			16'h2b9b: y = 16'h200;
			16'h2b9c: y = 16'h200;
			16'h2b9d: y = 16'h200;
			16'h2b9e: y = 16'h200;
			16'h2b9f: y = 16'h200;
			16'h2ba0: y = 16'h200;
			16'h2ba1: y = 16'h200;
			16'h2ba2: y = 16'h200;
			16'h2ba3: y = 16'h200;
			16'h2ba4: y = 16'h200;
			16'h2ba5: y = 16'h200;
			16'h2ba6: y = 16'h200;
			16'h2ba7: y = 16'h200;
			16'h2ba8: y = 16'h200;
			16'h2ba9: y = 16'h200;
			16'h2baa: y = 16'h200;
			16'h2bab: y = 16'h200;
			16'h2bac: y = 16'h200;
			16'h2bad: y = 16'h200;
			16'h2bae: y = 16'h200;
			16'h2baf: y = 16'h200;
			16'h2bb0: y = 16'h200;
			16'h2bb1: y = 16'h200;
			16'h2bb2: y = 16'h200;
			16'h2bb3: y = 16'h200;
			16'h2bb4: y = 16'h200;
			16'h2bb5: y = 16'h200;
			16'h2bb6: y = 16'h200;
			16'h2bb7: y = 16'h200;
			16'h2bb8: y = 16'h200;
			16'h2bb9: y = 16'h200;
			16'h2bba: y = 16'h200;
			16'h2bbb: y = 16'h200;
			16'h2bbc: y = 16'h200;
			16'h2bbd: y = 16'h200;
			16'h2bbe: y = 16'h200;
			16'h2bbf: y = 16'h200;
			16'h2bc0: y = 16'h200;
			16'h2bc1: y = 16'h200;
			16'h2bc2: y = 16'h200;
			16'h2bc3: y = 16'h200;
			16'h2bc4: y = 16'h200;
			16'h2bc5: y = 16'h200;
			16'h2bc6: y = 16'h200;
			16'h2bc7: y = 16'h200;
			16'h2bc8: y = 16'h200;
			16'h2bc9: y = 16'h200;
			16'h2bca: y = 16'h200;
			16'h2bcb: y = 16'h200;
			16'h2bcc: y = 16'h200;
			16'h2bcd: y = 16'h200;
			16'h2bce: y = 16'h200;
			16'h2bcf: y = 16'h200;
			16'h2bd0: y = 16'h200;
			16'h2bd1: y = 16'h200;
			16'h2bd2: y = 16'h200;
			16'h2bd3: y = 16'h200;
			16'h2bd4: y = 16'h200;
			16'h2bd5: y = 16'h200;
			16'h2bd6: y = 16'h200;
			16'h2bd7: y = 16'h200;
			16'h2bd8: y = 16'h200;
			16'h2bd9: y = 16'h200;
			16'h2bda: y = 16'h200;
			16'h2bdb: y = 16'h200;
			16'h2bdc: y = 16'h200;
			16'h2bdd: y = 16'h200;
			16'h2bde: y = 16'h200;
			16'h2bdf: y = 16'h200;
			16'h2be0: y = 16'h200;
			16'h2be1: y = 16'h200;
			16'h2be2: y = 16'h200;
			16'h2be3: y = 16'h200;
			16'h2be4: y = 16'h200;
			16'h2be5: y = 16'h200;
			16'h2be6: y = 16'h200;
			16'h2be7: y = 16'h200;
			16'h2be8: y = 16'h200;
			16'h2be9: y = 16'h200;
			16'h2bea: y = 16'h200;
			16'h2beb: y = 16'h200;
			16'h2bec: y = 16'h200;
			16'h2bed: y = 16'h200;
			16'h2bee: y = 16'h200;
			16'h2bef: y = 16'h200;
			16'h2bf0: y = 16'h200;
			16'h2bf1: y = 16'h200;
			16'h2bf2: y = 16'h200;
			16'h2bf3: y = 16'h200;
			16'h2bf4: y = 16'h200;
			16'h2bf5: y = 16'h200;
			16'h2bf6: y = 16'h200;
			16'h2bf7: y = 16'h200;
			16'h2bf8: y = 16'h200;
			16'h2bf9: y = 16'h200;
			16'h2bfa: y = 16'h200;
			16'h2bfb: y = 16'h200;
			16'h2bfc: y = 16'h200;
			16'h2bfd: y = 16'h200;
			16'h2bfe: y = 16'h200;
			16'h2bff: y = 16'h200;
			16'h2c00: y = 16'h200;
			16'h2c01: y = 16'h200;
			16'h2c02: y = 16'h200;
			16'h2c03: y = 16'h200;
			16'h2c04: y = 16'h200;
			16'h2c05: y = 16'h200;
			16'h2c06: y = 16'h200;
			16'h2c07: y = 16'h200;
			16'h2c08: y = 16'h200;
			16'h2c09: y = 16'h200;
			16'h2c0a: y = 16'h200;
			16'h2c0b: y = 16'h200;
			16'h2c0c: y = 16'h200;
			16'h2c0d: y = 16'h200;
			16'h2c0e: y = 16'h200;
			16'h2c0f: y = 16'h200;
			16'h2c10: y = 16'h200;
			16'h2c11: y = 16'h200;
			16'h2c12: y = 16'h200;
			16'h2c13: y = 16'h200;
			16'h2c14: y = 16'h200;
			16'h2c15: y = 16'h200;
			16'h2c16: y = 16'h200;
			16'h2c17: y = 16'h200;
			16'h2c18: y = 16'h200;
			16'h2c19: y = 16'h200;
			16'h2c1a: y = 16'h200;
			16'h2c1b: y = 16'h200;
			16'h2c1c: y = 16'h200;
			16'h2c1d: y = 16'h200;
			16'h2c1e: y = 16'h200;
			16'h2c1f: y = 16'h200;
			16'h2c20: y = 16'h200;
			16'h2c21: y = 16'h200;
			16'h2c22: y = 16'h200;
			16'h2c23: y = 16'h200;
			16'h2c24: y = 16'h200;
			16'h2c25: y = 16'h200;
			16'h2c26: y = 16'h200;
			16'h2c27: y = 16'h200;
			16'h2c28: y = 16'h200;
			16'h2c29: y = 16'h200;
			16'h2c2a: y = 16'h200;
			16'h2c2b: y = 16'h200;
			16'h2c2c: y = 16'h200;
			16'h2c2d: y = 16'h200;
			16'h2c2e: y = 16'h200;
			16'h2c2f: y = 16'h200;
			16'h2c30: y = 16'h200;
			16'h2c31: y = 16'h200;
			16'h2c32: y = 16'h200;
			16'h2c33: y = 16'h200;
			16'h2c34: y = 16'h200;
			16'h2c35: y = 16'h200;
			16'h2c36: y = 16'h200;
			16'h2c37: y = 16'h200;
			16'h2c38: y = 16'h200;
			16'h2c39: y = 16'h200;
			16'h2c3a: y = 16'h200;
			16'h2c3b: y = 16'h200;
			16'h2c3c: y = 16'h200;
			16'h2c3d: y = 16'h200;
			16'h2c3e: y = 16'h200;
			16'h2c3f: y = 16'h200;
			16'h2c40: y = 16'h200;
			16'h2c41: y = 16'h200;
			16'h2c42: y = 16'h200;
			16'h2c43: y = 16'h200;
			16'h2c44: y = 16'h200;
			16'h2c45: y = 16'h200;
			16'h2c46: y = 16'h200;
			16'h2c47: y = 16'h200;
			16'h2c48: y = 16'h200;
			16'h2c49: y = 16'h200;
			16'h2c4a: y = 16'h200;
			16'h2c4b: y = 16'h200;
			16'h2c4c: y = 16'h200;
			16'h2c4d: y = 16'h200;
			16'h2c4e: y = 16'h200;
			16'h2c4f: y = 16'h200;
			16'h2c50: y = 16'h200;
			16'h2c51: y = 16'h200;
			16'h2c52: y = 16'h200;
			16'h2c53: y = 16'h200;
			16'h2c54: y = 16'h200;
			16'h2c55: y = 16'h200;
			16'h2c56: y = 16'h200;
			16'h2c57: y = 16'h200;
			16'h2c58: y = 16'h200;
			16'h2c59: y = 16'h200;
			16'h2c5a: y = 16'h200;
			16'h2c5b: y = 16'h200;
			16'h2c5c: y = 16'h200;
			16'h2c5d: y = 16'h200;
			16'h2c5e: y = 16'h200;
			16'h2c5f: y = 16'h200;
			16'h2c60: y = 16'h200;
			16'h2c61: y = 16'h200;
			16'h2c62: y = 16'h200;
			16'h2c63: y = 16'h200;
			16'h2c64: y = 16'h200;
			16'h2c65: y = 16'h200;
			16'h2c66: y = 16'h200;
			16'h2c67: y = 16'h200;
			16'h2c68: y = 16'h200;
			16'h2c69: y = 16'h200;
			16'h2c6a: y = 16'h200;
			16'h2c6b: y = 16'h200;
			16'h2c6c: y = 16'h200;
			16'h2c6d: y = 16'h200;
			16'h2c6e: y = 16'h200;
			16'h2c6f: y = 16'h200;
			16'h2c70: y = 16'h200;
			16'h2c71: y = 16'h200;
			16'h2c72: y = 16'h200;
			16'h2c73: y = 16'h200;
			16'h2c74: y = 16'h200;
			16'h2c75: y = 16'h200;
			16'h2c76: y = 16'h200;
			16'h2c77: y = 16'h200;
			16'h2c78: y = 16'h200;
			16'h2c79: y = 16'h200;
			16'h2c7a: y = 16'h200;
			16'h2c7b: y = 16'h200;
			16'h2c7c: y = 16'h200;
			16'h2c7d: y = 16'h200;
			16'h2c7e: y = 16'h200;
			16'h2c7f: y = 16'h200;
			16'h2c80: y = 16'h200;
			16'h2c81: y = 16'h200;
			16'h2c82: y = 16'h200;
			16'h2c83: y = 16'h200;
			16'h2c84: y = 16'h200;
			16'h2c85: y = 16'h200;
			16'h2c86: y = 16'h200;
			16'h2c87: y = 16'h200;
			16'h2c88: y = 16'h200;
			16'h2c89: y = 16'h200;
			16'h2c8a: y = 16'h200;
			16'h2c8b: y = 16'h200;
			16'h2c8c: y = 16'h200;
			16'h2c8d: y = 16'h200;
			16'h2c8e: y = 16'h200;
			16'h2c8f: y = 16'h200;
			16'h2c90: y = 16'h200;
			16'h2c91: y = 16'h200;
			16'h2c92: y = 16'h200;
			16'h2c93: y = 16'h200;
			16'h2c94: y = 16'h200;
			16'h2c95: y = 16'h200;
			16'h2c96: y = 16'h200;
			16'h2c97: y = 16'h200;
			16'h2c98: y = 16'h200;
			16'h2c99: y = 16'h200;
			16'h2c9a: y = 16'h200;
			16'h2c9b: y = 16'h200;
			16'h2c9c: y = 16'h200;
			16'h2c9d: y = 16'h200;
			16'h2c9e: y = 16'h200;
			16'h2c9f: y = 16'h200;
			16'h2ca0: y = 16'h200;
			16'h2ca1: y = 16'h200;
			16'h2ca2: y = 16'h200;
			16'h2ca3: y = 16'h200;
			16'h2ca4: y = 16'h200;
			16'h2ca5: y = 16'h200;
			16'h2ca6: y = 16'h200;
			16'h2ca7: y = 16'h200;
			16'h2ca8: y = 16'h200;
			16'h2ca9: y = 16'h200;
			16'h2caa: y = 16'h200;
			16'h2cab: y = 16'h200;
			16'h2cac: y = 16'h200;
			16'h2cad: y = 16'h200;
			16'h2cae: y = 16'h200;
			16'h2caf: y = 16'h200;
			16'h2cb0: y = 16'h200;
			16'h2cb1: y = 16'h200;
			16'h2cb2: y = 16'h200;
			16'h2cb3: y = 16'h200;
			16'h2cb4: y = 16'h200;
			16'h2cb5: y = 16'h200;
			16'h2cb6: y = 16'h200;
			16'h2cb7: y = 16'h200;
			16'h2cb8: y = 16'h200;
			16'h2cb9: y = 16'h200;
			16'h2cba: y = 16'h200;
			16'h2cbb: y = 16'h200;
			16'h2cbc: y = 16'h200;
			16'h2cbd: y = 16'h200;
			16'h2cbe: y = 16'h200;
			16'h2cbf: y = 16'h200;
			16'h2cc0: y = 16'h200;
			16'h2cc1: y = 16'h200;
			16'h2cc2: y = 16'h200;
			16'h2cc3: y = 16'h200;
			16'h2cc4: y = 16'h200;
			16'h2cc5: y = 16'h200;
			16'h2cc6: y = 16'h200;
			16'h2cc7: y = 16'h200;
			16'h2cc8: y = 16'h200;
			16'h2cc9: y = 16'h200;
			16'h2cca: y = 16'h200;
			16'h2ccb: y = 16'h200;
			16'h2ccc: y = 16'h200;
			16'h2ccd: y = 16'h200;
			16'h2cce: y = 16'h200;
			16'h2ccf: y = 16'h200;
			16'h2cd0: y = 16'h200;
			16'h2cd1: y = 16'h200;
			16'h2cd2: y = 16'h200;
			16'h2cd3: y = 16'h200;
			16'h2cd4: y = 16'h200;
			16'h2cd5: y = 16'h200;
			16'h2cd6: y = 16'h200;
			16'h2cd7: y = 16'h200;
			16'h2cd8: y = 16'h200;
			16'h2cd9: y = 16'h200;
			16'h2cda: y = 16'h200;
			16'h2cdb: y = 16'h200;
			16'h2cdc: y = 16'h200;
			16'h2cdd: y = 16'h200;
			16'h2cde: y = 16'h200;
			16'h2cdf: y = 16'h200;
			16'h2ce0: y = 16'h200;
			16'h2ce1: y = 16'h200;
			16'h2ce2: y = 16'h200;
			16'h2ce3: y = 16'h200;
			16'h2ce4: y = 16'h200;
			16'h2ce5: y = 16'h200;
			16'h2ce6: y = 16'h200;
			16'h2ce7: y = 16'h200;
			16'h2ce8: y = 16'h200;
			16'h2ce9: y = 16'h200;
			16'h2cea: y = 16'h200;
			16'h2ceb: y = 16'h200;
			16'h2cec: y = 16'h200;
			16'h2ced: y = 16'h200;
			16'h2cee: y = 16'h200;
			16'h2cef: y = 16'h200;
			16'h2cf0: y = 16'h200;
			16'h2cf1: y = 16'h200;
			16'h2cf2: y = 16'h200;
			16'h2cf3: y = 16'h200;
			16'h2cf4: y = 16'h200;
			16'h2cf5: y = 16'h200;
			16'h2cf6: y = 16'h200;
			16'h2cf7: y = 16'h200;
			16'h2cf8: y = 16'h200;
			16'h2cf9: y = 16'h200;
			16'h2cfa: y = 16'h200;
			16'h2cfb: y = 16'h200;
			16'h2cfc: y = 16'h200;
			16'h2cfd: y = 16'h200;
			16'h2cfe: y = 16'h200;
			16'h2cff: y = 16'h200;
			16'h2d00: y = 16'h200;
			16'h2d01: y = 16'h200;
			16'h2d02: y = 16'h200;
			16'h2d03: y = 16'h200;
			16'h2d04: y = 16'h200;
			16'h2d05: y = 16'h200;
			16'h2d06: y = 16'h200;
			16'h2d07: y = 16'h200;
			16'h2d08: y = 16'h200;
			16'h2d09: y = 16'h200;
			16'h2d0a: y = 16'h200;
			16'h2d0b: y = 16'h200;
			16'h2d0c: y = 16'h200;
			16'h2d0d: y = 16'h200;
			16'h2d0e: y = 16'h200;
			16'h2d0f: y = 16'h200;
			16'h2d10: y = 16'h200;
			16'h2d11: y = 16'h200;
			16'h2d12: y = 16'h200;
			16'h2d13: y = 16'h200;
			16'h2d14: y = 16'h200;
			16'h2d15: y = 16'h200;
			16'h2d16: y = 16'h200;
			16'h2d17: y = 16'h200;
			16'h2d18: y = 16'h200;
			16'h2d19: y = 16'h200;
			16'h2d1a: y = 16'h200;
			16'h2d1b: y = 16'h200;
			16'h2d1c: y = 16'h200;
			16'h2d1d: y = 16'h200;
			16'h2d1e: y = 16'h200;
			16'h2d1f: y = 16'h200;
			16'h2d20: y = 16'h200;
			16'h2d21: y = 16'h200;
			16'h2d22: y = 16'h200;
			16'h2d23: y = 16'h200;
			16'h2d24: y = 16'h200;
			16'h2d25: y = 16'h200;
			16'h2d26: y = 16'h200;
			16'h2d27: y = 16'h200;
			16'h2d28: y = 16'h200;
			16'h2d29: y = 16'h200;
			16'h2d2a: y = 16'h200;
			16'h2d2b: y = 16'h200;
			16'h2d2c: y = 16'h200;
			16'h2d2d: y = 16'h200;
			16'h2d2e: y = 16'h200;
			16'h2d2f: y = 16'h200;
			16'h2d30: y = 16'h200;
			16'h2d31: y = 16'h200;
			16'h2d32: y = 16'h200;
			16'h2d33: y = 16'h200;
			16'h2d34: y = 16'h200;
			16'h2d35: y = 16'h200;
			16'h2d36: y = 16'h200;
			16'h2d37: y = 16'h200;
			16'h2d38: y = 16'h200;
			16'h2d39: y = 16'h200;
			16'h2d3a: y = 16'h200;
			16'h2d3b: y = 16'h200;
			16'h2d3c: y = 16'h200;
			16'h2d3d: y = 16'h200;
			16'h2d3e: y = 16'h200;
			16'h2d3f: y = 16'h200;
			16'h2d40: y = 16'h200;
			16'h2d41: y = 16'h200;
			16'h2d42: y = 16'h200;
			16'h2d43: y = 16'h200;
			16'h2d44: y = 16'h200;
			16'h2d45: y = 16'h200;
			16'h2d46: y = 16'h200;
			16'h2d47: y = 16'h200;
			16'h2d48: y = 16'h200;
			16'h2d49: y = 16'h200;
			16'h2d4a: y = 16'h200;
			16'h2d4b: y = 16'h200;
			16'h2d4c: y = 16'h200;
			16'h2d4d: y = 16'h200;
			16'h2d4e: y = 16'h200;
			16'h2d4f: y = 16'h200;
			16'h2d50: y = 16'h200;
			16'h2d51: y = 16'h200;
			16'h2d52: y = 16'h200;
			16'h2d53: y = 16'h200;
			16'h2d54: y = 16'h200;
			16'h2d55: y = 16'h200;
			16'h2d56: y = 16'h200;
			16'h2d57: y = 16'h200;
			16'h2d58: y = 16'h200;
			16'h2d59: y = 16'h200;
			16'h2d5a: y = 16'h200;
			16'h2d5b: y = 16'h200;
			16'h2d5c: y = 16'h200;
			16'h2d5d: y = 16'h200;
			16'h2d5e: y = 16'h200;
			16'h2d5f: y = 16'h200;
			16'h2d60: y = 16'h200;
			16'h2d61: y = 16'h200;
			16'h2d62: y = 16'h200;
			16'h2d63: y = 16'h200;
			16'h2d64: y = 16'h200;
			16'h2d65: y = 16'h200;
			16'h2d66: y = 16'h200;
			16'h2d67: y = 16'h200;
			16'h2d68: y = 16'h200;
			16'h2d69: y = 16'h200;
			16'h2d6a: y = 16'h200;
			16'h2d6b: y = 16'h200;
			16'h2d6c: y = 16'h200;
			16'h2d6d: y = 16'h200;
			16'h2d6e: y = 16'h200;
			16'h2d6f: y = 16'h200;
			16'h2d70: y = 16'h200;
			16'h2d71: y = 16'h200;
			16'h2d72: y = 16'h200;
			16'h2d73: y = 16'h200;
			16'h2d74: y = 16'h200;
			16'h2d75: y = 16'h200;
			16'h2d76: y = 16'h200;
			16'h2d77: y = 16'h200;
			16'h2d78: y = 16'h200;
			16'h2d79: y = 16'h200;
			16'h2d7a: y = 16'h200;
			16'h2d7b: y = 16'h200;
			16'h2d7c: y = 16'h200;
			16'h2d7d: y = 16'h200;
			16'h2d7e: y = 16'h200;
			16'h2d7f: y = 16'h200;
			16'h2d80: y = 16'h200;
			16'h2d81: y = 16'h200;
			16'h2d82: y = 16'h200;
			16'h2d83: y = 16'h200;
			16'h2d84: y = 16'h200;
			16'h2d85: y = 16'h200;
			16'h2d86: y = 16'h200;
			16'h2d87: y = 16'h200;
			16'h2d88: y = 16'h200;
			16'h2d89: y = 16'h200;
			16'h2d8a: y = 16'h200;
			16'h2d8b: y = 16'h200;
			16'h2d8c: y = 16'h200;
			16'h2d8d: y = 16'h200;
			16'h2d8e: y = 16'h200;
			16'h2d8f: y = 16'h200;
			16'h2d90: y = 16'h200;
			16'h2d91: y = 16'h200;
			16'h2d92: y = 16'h200;
			16'h2d93: y = 16'h200;
			16'h2d94: y = 16'h200;
			16'h2d95: y = 16'h200;
			16'h2d96: y = 16'h200;
			16'h2d97: y = 16'h200;
			16'h2d98: y = 16'h200;
			16'h2d99: y = 16'h200;
			16'h2d9a: y = 16'h200;
			16'h2d9b: y = 16'h200;
			16'h2d9c: y = 16'h200;
			16'h2d9d: y = 16'h200;
			16'h2d9e: y = 16'h200;
			16'h2d9f: y = 16'h200;
			16'h2da0: y = 16'h200;
			16'h2da1: y = 16'h200;
			16'h2da2: y = 16'h200;
			16'h2da3: y = 16'h200;
			16'h2da4: y = 16'h200;
			16'h2da5: y = 16'h200;
			16'h2da6: y = 16'h200;
			16'h2da7: y = 16'h200;
			16'h2da8: y = 16'h200;
			16'h2da9: y = 16'h200;
			16'h2daa: y = 16'h200;
			16'h2dab: y = 16'h200;
			16'h2dac: y = 16'h200;
			16'h2dad: y = 16'h200;
			16'h2dae: y = 16'h200;
			16'h2daf: y = 16'h200;
			16'h2db0: y = 16'h200;
			16'h2db1: y = 16'h200;
			16'h2db2: y = 16'h200;
			16'h2db3: y = 16'h200;
			16'h2db4: y = 16'h200;
			16'h2db5: y = 16'h200;
			16'h2db6: y = 16'h200;
			16'h2db7: y = 16'h200;
			16'h2db8: y = 16'h200;
			16'h2db9: y = 16'h200;
			16'h2dba: y = 16'h200;
			16'h2dbb: y = 16'h200;
			16'h2dbc: y = 16'h200;
			16'h2dbd: y = 16'h200;
			16'h2dbe: y = 16'h200;
			16'h2dbf: y = 16'h200;
			16'h2dc0: y = 16'h200;
			16'h2dc1: y = 16'h200;
			16'h2dc2: y = 16'h200;
			16'h2dc3: y = 16'h200;
			16'h2dc4: y = 16'h200;
			16'h2dc5: y = 16'h200;
			16'h2dc6: y = 16'h200;
			16'h2dc7: y = 16'h200;
			16'h2dc8: y = 16'h200;
			16'h2dc9: y = 16'h200;
			16'h2dca: y = 16'h200;
			16'h2dcb: y = 16'h200;
			16'h2dcc: y = 16'h200;
			16'h2dcd: y = 16'h200;
			16'h2dce: y = 16'h200;
			16'h2dcf: y = 16'h200;
			16'h2dd0: y = 16'h200;
			16'h2dd1: y = 16'h200;
			16'h2dd2: y = 16'h200;
			16'h2dd3: y = 16'h200;
			16'h2dd4: y = 16'h200;
			16'h2dd5: y = 16'h200;
			16'h2dd6: y = 16'h200;
			16'h2dd7: y = 16'h200;
			16'h2dd8: y = 16'h200;
			16'h2dd9: y = 16'h200;
			16'h2dda: y = 16'h200;
			16'h2ddb: y = 16'h200;
			16'h2ddc: y = 16'h200;
			16'h2ddd: y = 16'h200;
			16'h2dde: y = 16'h200;
			16'h2ddf: y = 16'h200;
			16'h2de0: y = 16'h200;
			16'h2de1: y = 16'h200;
			16'h2de2: y = 16'h200;
			16'h2de3: y = 16'h200;
			16'h2de4: y = 16'h200;
			16'h2de5: y = 16'h200;
			16'h2de6: y = 16'h200;
			16'h2de7: y = 16'h200;
			16'h2de8: y = 16'h200;
			16'h2de9: y = 16'h200;
			16'h2dea: y = 16'h200;
			16'h2deb: y = 16'h200;
			16'h2dec: y = 16'h200;
			16'h2ded: y = 16'h200;
			16'h2dee: y = 16'h200;
			16'h2def: y = 16'h200;
			16'h2df0: y = 16'h200;
			16'h2df1: y = 16'h200;
			16'h2df2: y = 16'h200;
			16'h2df3: y = 16'h200;
			16'h2df4: y = 16'h200;
			16'h2df5: y = 16'h200;
			16'h2df6: y = 16'h200;
			16'h2df7: y = 16'h200;
			16'h2df8: y = 16'h200;
			16'h2df9: y = 16'h200;
			16'h2dfa: y = 16'h200;
			16'h2dfb: y = 16'h200;
			16'h2dfc: y = 16'h200;
			16'h2dfd: y = 16'h200;
			16'h2dfe: y = 16'h200;
			16'h2dff: y = 16'h200;
			16'h2e00: y = 16'h200;
			16'h2e01: y = 16'h200;
			16'h2e02: y = 16'h200;
			16'h2e03: y = 16'h200;
			16'h2e04: y = 16'h200;
			16'h2e05: y = 16'h200;
			16'h2e06: y = 16'h200;
			16'h2e07: y = 16'h200;
			16'h2e08: y = 16'h200;
			16'h2e09: y = 16'h200;
			16'h2e0a: y = 16'h200;
			16'h2e0b: y = 16'h200;
			16'h2e0c: y = 16'h200;
			16'h2e0d: y = 16'h200;
			16'h2e0e: y = 16'h200;
			16'h2e0f: y = 16'h200;
			16'h2e10: y = 16'h200;
			16'h2e11: y = 16'h200;
			16'h2e12: y = 16'h200;
			16'h2e13: y = 16'h200;
			16'h2e14: y = 16'h200;
			16'h2e15: y = 16'h200;
			16'h2e16: y = 16'h200;
			16'h2e17: y = 16'h200;
			16'h2e18: y = 16'h200;
			16'h2e19: y = 16'h200;
			16'h2e1a: y = 16'h200;
			16'h2e1b: y = 16'h200;
			16'h2e1c: y = 16'h200;
			16'h2e1d: y = 16'h200;
			16'h2e1e: y = 16'h200;
			16'h2e1f: y = 16'h200;
			16'h2e20: y = 16'h200;
			16'h2e21: y = 16'h200;
			16'h2e22: y = 16'h200;
			16'h2e23: y = 16'h200;
			16'h2e24: y = 16'h200;
			16'h2e25: y = 16'h200;
			16'h2e26: y = 16'h200;
			16'h2e27: y = 16'h200;
			16'h2e28: y = 16'h200;
			16'h2e29: y = 16'h200;
			16'h2e2a: y = 16'h200;
			16'h2e2b: y = 16'h200;
			16'h2e2c: y = 16'h200;
			16'h2e2d: y = 16'h200;
			16'h2e2e: y = 16'h200;
			16'h2e2f: y = 16'h200;
			16'h2e30: y = 16'h200;
			16'h2e31: y = 16'h200;
			16'h2e32: y = 16'h200;
			16'h2e33: y = 16'h200;
			16'h2e34: y = 16'h200;
			16'h2e35: y = 16'h200;
			16'h2e36: y = 16'h200;
			16'h2e37: y = 16'h200;
			16'h2e38: y = 16'h200;
			16'h2e39: y = 16'h200;
			16'h2e3a: y = 16'h200;
			16'h2e3b: y = 16'h200;
			16'h2e3c: y = 16'h200;
			16'h2e3d: y = 16'h200;
			16'h2e3e: y = 16'h200;
			16'h2e3f: y = 16'h200;
			16'h2e40: y = 16'h200;
			16'h2e41: y = 16'h200;
			16'h2e42: y = 16'h200;
			16'h2e43: y = 16'h200;
			16'h2e44: y = 16'h200;
			16'h2e45: y = 16'h200;
			16'h2e46: y = 16'h200;
			16'h2e47: y = 16'h200;
			16'h2e48: y = 16'h200;
			16'h2e49: y = 16'h200;
			16'h2e4a: y = 16'h200;
			16'h2e4b: y = 16'h200;
			16'h2e4c: y = 16'h200;
			16'h2e4d: y = 16'h200;
			16'h2e4e: y = 16'h200;
			16'h2e4f: y = 16'h200;
			16'h2e50: y = 16'h200;
			16'h2e51: y = 16'h200;
			16'h2e52: y = 16'h200;
			16'h2e53: y = 16'h200;
			16'h2e54: y = 16'h200;
			16'h2e55: y = 16'h200;
			16'h2e56: y = 16'h200;
			16'h2e57: y = 16'h200;
			16'h2e58: y = 16'h200;
			16'h2e59: y = 16'h200;
			16'h2e5a: y = 16'h200;
			16'h2e5b: y = 16'h200;
			16'h2e5c: y = 16'h200;
			16'h2e5d: y = 16'h200;
			16'h2e5e: y = 16'h200;
			16'h2e5f: y = 16'h200;
			16'h2e60: y = 16'h200;
			16'h2e61: y = 16'h200;
			16'h2e62: y = 16'h200;
			16'h2e63: y = 16'h200;
			16'h2e64: y = 16'h200;
			16'h2e65: y = 16'h200;
			16'h2e66: y = 16'h200;
			16'h2e67: y = 16'h200;
			16'h2e68: y = 16'h200;
			16'h2e69: y = 16'h200;
			16'h2e6a: y = 16'h200;
			16'h2e6b: y = 16'h200;
			16'h2e6c: y = 16'h200;
			16'h2e6d: y = 16'h200;
			16'h2e6e: y = 16'h200;
			16'h2e6f: y = 16'h200;
			16'h2e70: y = 16'h200;
			16'h2e71: y = 16'h200;
			16'h2e72: y = 16'h200;
			16'h2e73: y = 16'h200;
			16'h2e74: y = 16'h200;
			16'h2e75: y = 16'h200;
			16'h2e76: y = 16'h200;
			16'h2e77: y = 16'h200;
			16'h2e78: y = 16'h200;
			16'h2e79: y = 16'h200;
			16'h2e7a: y = 16'h200;
			16'h2e7b: y = 16'h200;
			16'h2e7c: y = 16'h200;
			16'h2e7d: y = 16'h200;
			16'h2e7e: y = 16'h200;
			16'h2e7f: y = 16'h200;
			16'h2e80: y = 16'h200;
			16'h2e81: y = 16'h200;
			16'h2e82: y = 16'h200;
			16'h2e83: y = 16'h200;
			16'h2e84: y = 16'h200;
			16'h2e85: y = 16'h200;
			16'h2e86: y = 16'h200;
			16'h2e87: y = 16'h200;
			16'h2e88: y = 16'h200;
			16'h2e89: y = 16'h200;
			16'h2e8a: y = 16'h200;
			16'h2e8b: y = 16'h200;
			16'h2e8c: y = 16'h200;
			16'h2e8d: y = 16'h200;
			16'h2e8e: y = 16'h200;
			16'h2e8f: y = 16'h200;
			16'h2e90: y = 16'h200;
			16'h2e91: y = 16'h200;
			16'h2e92: y = 16'h200;
			16'h2e93: y = 16'h200;
			16'h2e94: y = 16'h200;
			16'h2e95: y = 16'h200;
			16'h2e96: y = 16'h200;
			16'h2e97: y = 16'h200;
			16'h2e98: y = 16'h200;
			16'h2e99: y = 16'h200;
			16'h2e9a: y = 16'h200;
			16'h2e9b: y = 16'h200;
			16'h2e9c: y = 16'h200;
			16'h2e9d: y = 16'h200;
			16'h2e9e: y = 16'h200;
			16'h2e9f: y = 16'h200;
			16'h2ea0: y = 16'h200;
			16'h2ea1: y = 16'h200;
			16'h2ea2: y = 16'h200;
			16'h2ea3: y = 16'h200;
			16'h2ea4: y = 16'h200;
			16'h2ea5: y = 16'h200;
			16'h2ea6: y = 16'h200;
			16'h2ea7: y = 16'h200;
			16'h2ea8: y = 16'h200;
			16'h2ea9: y = 16'h200;
			16'h2eaa: y = 16'h200;
			16'h2eab: y = 16'h200;
			16'h2eac: y = 16'h200;
			16'h2ead: y = 16'h200;
			16'h2eae: y = 16'h200;
			16'h2eaf: y = 16'h200;
			16'h2eb0: y = 16'h200;
			16'h2eb1: y = 16'h200;
			16'h2eb2: y = 16'h200;
			16'h2eb3: y = 16'h200;
			16'h2eb4: y = 16'h200;
			16'h2eb5: y = 16'h200;
			16'h2eb6: y = 16'h200;
			16'h2eb7: y = 16'h200;
			16'h2eb8: y = 16'h200;
			16'h2eb9: y = 16'h200;
			16'h2eba: y = 16'h200;
			16'h2ebb: y = 16'h200;
			16'h2ebc: y = 16'h200;
			16'h2ebd: y = 16'h200;
			16'h2ebe: y = 16'h200;
			16'h2ebf: y = 16'h200;
			16'h2ec0: y = 16'h200;
			16'h2ec1: y = 16'h200;
			16'h2ec2: y = 16'h200;
			16'h2ec3: y = 16'h200;
			16'h2ec4: y = 16'h200;
			16'h2ec5: y = 16'h200;
			16'h2ec6: y = 16'h200;
			16'h2ec7: y = 16'h200;
			16'h2ec8: y = 16'h200;
			16'h2ec9: y = 16'h200;
			16'h2eca: y = 16'h200;
			16'h2ecb: y = 16'h200;
			16'h2ecc: y = 16'h200;
			16'h2ecd: y = 16'h200;
			16'h2ece: y = 16'h200;
			16'h2ecf: y = 16'h200;
			16'h2ed0: y = 16'h200;
			16'h2ed1: y = 16'h200;
			16'h2ed2: y = 16'h200;
			16'h2ed3: y = 16'h200;
			16'h2ed4: y = 16'h200;
			16'h2ed5: y = 16'h200;
			16'h2ed6: y = 16'h200;
			16'h2ed7: y = 16'h200;
			16'h2ed8: y = 16'h200;
			16'h2ed9: y = 16'h200;
			16'h2eda: y = 16'h200;
			16'h2edb: y = 16'h200;
			16'h2edc: y = 16'h200;
			16'h2edd: y = 16'h200;
			16'h2ede: y = 16'h200;
			16'h2edf: y = 16'h200;
			16'h2ee0: y = 16'h200;
			16'h2ee1: y = 16'h200;
			16'h2ee2: y = 16'h200;
			16'h2ee3: y = 16'h200;
			16'h2ee4: y = 16'h200;
			16'h2ee5: y = 16'h200;
			16'h2ee6: y = 16'h200;
			16'h2ee7: y = 16'h200;
			16'h2ee8: y = 16'h200;
			16'h2ee9: y = 16'h200;
			16'h2eea: y = 16'h200;
			16'h2eeb: y = 16'h200;
			16'h2eec: y = 16'h200;
			16'h2eed: y = 16'h200;
			16'h2eee: y = 16'h200;
			16'h2eef: y = 16'h200;
			16'h2ef0: y = 16'h200;
			16'h2ef1: y = 16'h200;
			16'h2ef2: y = 16'h200;
			16'h2ef3: y = 16'h200;
			16'h2ef4: y = 16'h200;
			16'h2ef5: y = 16'h200;
			16'h2ef6: y = 16'h200;
			16'h2ef7: y = 16'h200;
			16'h2ef8: y = 16'h200;
			16'h2ef9: y = 16'h200;
			16'h2efa: y = 16'h200;
			16'h2efb: y = 16'h200;
			16'h2efc: y = 16'h200;
			16'h2efd: y = 16'h200;
			16'h2efe: y = 16'h200;
			16'h2eff: y = 16'h200;
			16'h2f00: y = 16'h200;
			16'h2f01: y = 16'h200;
			16'h2f02: y = 16'h200;
			16'h2f03: y = 16'h200;
			16'h2f04: y = 16'h200;
			16'h2f05: y = 16'h200;
			16'h2f06: y = 16'h200;
			16'h2f07: y = 16'h200;
			16'h2f08: y = 16'h200;
			16'h2f09: y = 16'h200;
			16'h2f0a: y = 16'h200;
			16'h2f0b: y = 16'h200;
			16'h2f0c: y = 16'h200;
			16'h2f0d: y = 16'h200;
			16'h2f0e: y = 16'h200;
			16'h2f0f: y = 16'h200;
			16'h2f10: y = 16'h200;
			16'h2f11: y = 16'h200;
			16'h2f12: y = 16'h200;
			16'h2f13: y = 16'h200;
			16'h2f14: y = 16'h200;
			16'h2f15: y = 16'h200;
			16'h2f16: y = 16'h200;
			16'h2f17: y = 16'h200;
			16'h2f18: y = 16'h200;
			16'h2f19: y = 16'h200;
			16'h2f1a: y = 16'h200;
			16'h2f1b: y = 16'h200;
			16'h2f1c: y = 16'h200;
			16'h2f1d: y = 16'h200;
			16'h2f1e: y = 16'h200;
			16'h2f1f: y = 16'h200;
			16'h2f20: y = 16'h200;
			16'h2f21: y = 16'h200;
			16'h2f22: y = 16'h200;
			16'h2f23: y = 16'h200;
			16'h2f24: y = 16'h200;
			16'h2f25: y = 16'h200;
			16'h2f26: y = 16'h200;
			16'h2f27: y = 16'h200;
			16'h2f28: y = 16'h200;
			16'h2f29: y = 16'h200;
			16'h2f2a: y = 16'h200;
			16'h2f2b: y = 16'h200;
			16'h2f2c: y = 16'h200;
			16'h2f2d: y = 16'h200;
			16'h2f2e: y = 16'h200;
			16'h2f2f: y = 16'h200;
			16'h2f30: y = 16'h200;
			16'h2f31: y = 16'h200;
			16'h2f32: y = 16'h200;
			16'h2f33: y = 16'h200;
			16'h2f34: y = 16'h200;
			16'h2f35: y = 16'h200;
			16'h2f36: y = 16'h200;
			16'h2f37: y = 16'h200;
			16'h2f38: y = 16'h200;
			16'h2f39: y = 16'h200;
			16'h2f3a: y = 16'h200;
			16'h2f3b: y = 16'h200;
			16'h2f3c: y = 16'h200;
			16'h2f3d: y = 16'h200;
			16'h2f3e: y = 16'h200;
			16'h2f3f: y = 16'h200;
			16'h2f40: y = 16'h200;
			16'h2f41: y = 16'h200;
			16'h2f42: y = 16'h200;
			16'h2f43: y = 16'h200;
			16'h2f44: y = 16'h200;
			16'h2f45: y = 16'h200;
			16'h2f46: y = 16'h200;
			16'h2f47: y = 16'h200;
			16'h2f48: y = 16'h200;
			16'h2f49: y = 16'h200;
			16'h2f4a: y = 16'h200;
			16'h2f4b: y = 16'h200;
			16'h2f4c: y = 16'h200;
			16'h2f4d: y = 16'h200;
			16'h2f4e: y = 16'h200;
			16'h2f4f: y = 16'h200;
			16'h2f50: y = 16'h200;
			16'h2f51: y = 16'h200;
			16'h2f52: y = 16'h200;
			16'h2f53: y = 16'h200;
			16'h2f54: y = 16'h200;
			16'h2f55: y = 16'h200;
			16'h2f56: y = 16'h200;
			16'h2f57: y = 16'h200;
			16'h2f58: y = 16'h200;
			16'h2f59: y = 16'h200;
			16'h2f5a: y = 16'h200;
			16'h2f5b: y = 16'h200;
			16'h2f5c: y = 16'h200;
			16'h2f5d: y = 16'h200;
			16'h2f5e: y = 16'h200;
			16'h2f5f: y = 16'h200;
			16'h2f60: y = 16'h200;
			16'h2f61: y = 16'h200;
			16'h2f62: y = 16'h200;
			16'h2f63: y = 16'h200;
			16'h2f64: y = 16'h200;
			16'h2f65: y = 16'h200;
			16'h2f66: y = 16'h200;
			16'h2f67: y = 16'h200;
			16'h2f68: y = 16'h200;
			16'h2f69: y = 16'h200;
			16'h2f6a: y = 16'h200;
			16'h2f6b: y = 16'h200;
			16'h2f6c: y = 16'h200;
			16'h2f6d: y = 16'h200;
			16'h2f6e: y = 16'h200;
			16'h2f6f: y = 16'h200;
			16'h2f70: y = 16'h200;
			16'h2f71: y = 16'h200;
			16'h2f72: y = 16'h200;
			16'h2f73: y = 16'h200;
			16'h2f74: y = 16'h200;
			16'h2f75: y = 16'h200;
			16'h2f76: y = 16'h200;
			16'h2f77: y = 16'h200;
			16'h2f78: y = 16'h200;
			16'h2f79: y = 16'h200;
			16'h2f7a: y = 16'h200;
			16'h2f7b: y = 16'h200;
			16'h2f7c: y = 16'h200;
			16'h2f7d: y = 16'h200;
			16'h2f7e: y = 16'h200;
			16'h2f7f: y = 16'h200;
			16'h2f80: y = 16'h200;
			16'h2f81: y = 16'h200;
			16'h2f82: y = 16'h200;
			16'h2f83: y = 16'h200;
			16'h2f84: y = 16'h200;
			16'h2f85: y = 16'h200;
			16'h2f86: y = 16'h200;
			16'h2f87: y = 16'h200;
			16'h2f88: y = 16'h200;
			16'h2f89: y = 16'h200;
			16'h2f8a: y = 16'h200;
			16'h2f8b: y = 16'h200;
			16'h2f8c: y = 16'h200;
			16'h2f8d: y = 16'h200;
			16'h2f8e: y = 16'h200;
			16'h2f8f: y = 16'h200;
			16'h2f90: y = 16'h200;
			16'h2f91: y = 16'h200;
			16'h2f92: y = 16'h200;
			16'h2f93: y = 16'h200;
			16'h2f94: y = 16'h200;
			16'h2f95: y = 16'h200;
			16'h2f96: y = 16'h200;
			16'h2f97: y = 16'h200;
			16'h2f98: y = 16'h200;
			16'h2f99: y = 16'h200;
			16'h2f9a: y = 16'h200;
			16'h2f9b: y = 16'h200;
			16'h2f9c: y = 16'h200;
			16'h2f9d: y = 16'h200;
			16'h2f9e: y = 16'h200;
			16'h2f9f: y = 16'h200;
			16'h2fa0: y = 16'h200;
			16'h2fa1: y = 16'h200;
			16'h2fa2: y = 16'h200;
			16'h2fa3: y = 16'h200;
			16'h2fa4: y = 16'h200;
			16'h2fa5: y = 16'h200;
			16'h2fa6: y = 16'h200;
			16'h2fa7: y = 16'h200;
			16'h2fa8: y = 16'h200;
			16'h2fa9: y = 16'h200;
			16'h2faa: y = 16'h200;
			16'h2fab: y = 16'h200;
			16'h2fac: y = 16'h200;
			16'h2fad: y = 16'h200;
			16'h2fae: y = 16'h200;
			16'h2faf: y = 16'h200;
			16'h2fb0: y = 16'h200;
			16'h2fb1: y = 16'h200;
			16'h2fb2: y = 16'h200;
			16'h2fb3: y = 16'h200;
			16'h2fb4: y = 16'h200;
			16'h2fb5: y = 16'h200;
			16'h2fb6: y = 16'h200;
			16'h2fb7: y = 16'h200;
			16'h2fb8: y = 16'h200;
			16'h2fb9: y = 16'h200;
			16'h2fba: y = 16'h200;
			16'h2fbb: y = 16'h200;
			16'h2fbc: y = 16'h200;
			16'h2fbd: y = 16'h200;
			16'h2fbe: y = 16'h200;
			16'h2fbf: y = 16'h200;
			16'h2fc0: y = 16'h200;
			16'h2fc1: y = 16'h200;
			16'h2fc2: y = 16'h200;
			16'h2fc3: y = 16'h200;
			16'h2fc4: y = 16'h200;
			16'h2fc5: y = 16'h200;
			16'h2fc6: y = 16'h200;
			16'h2fc7: y = 16'h200;
			16'h2fc8: y = 16'h200;
			16'h2fc9: y = 16'h200;
			16'h2fca: y = 16'h200;
			16'h2fcb: y = 16'h200;
			16'h2fcc: y = 16'h200;
			16'h2fcd: y = 16'h200;
			16'h2fce: y = 16'h200;
			16'h2fcf: y = 16'h200;
			16'h2fd0: y = 16'h200;
			16'h2fd1: y = 16'h200;
			16'h2fd2: y = 16'h200;
			16'h2fd3: y = 16'h200;
			16'h2fd4: y = 16'h200;
			16'h2fd5: y = 16'h200;
			16'h2fd6: y = 16'h200;
			16'h2fd7: y = 16'h200;
			16'h2fd8: y = 16'h200;
			16'h2fd9: y = 16'h200;
			16'h2fda: y = 16'h200;
			16'h2fdb: y = 16'h200;
			16'h2fdc: y = 16'h200;
			16'h2fdd: y = 16'h200;
			16'h2fde: y = 16'h200;
			16'h2fdf: y = 16'h200;
			16'h2fe0: y = 16'h200;
			16'h2fe1: y = 16'h200;
			16'h2fe2: y = 16'h200;
			16'h2fe3: y = 16'h200;
			16'h2fe4: y = 16'h200;
			16'h2fe5: y = 16'h200;
			16'h2fe6: y = 16'h200;
			16'h2fe7: y = 16'h200;
			16'h2fe8: y = 16'h200;
			16'h2fe9: y = 16'h200;
			16'h2fea: y = 16'h200;
			16'h2feb: y = 16'h200;
			16'h2fec: y = 16'h200;
			16'h2fed: y = 16'h200;
			16'h2fee: y = 16'h200;
			16'h2fef: y = 16'h200;
			16'h2ff0: y = 16'h200;
			16'h2ff1: y = 16'h200;
			16'h2ff2: y = 16'h200;
			16'h2ff3: y = 16'h200;
			16'h2ff4: y = 16'h200;
			16'h2ff5: y = 16'h200;
			16'h2ff6: y = 16'h200;
			16'h2ff7: y = 16'h200;
			16'h2ff8: y = 16'h200;
			16'h2ff9: y = 16'h200;
			16'h2ffa: y = 16'h200;
			16'h2ffb: y = 16'h200;
			16'h2ffc: y = 16'h200;
			16'h2ffd: y = 16'h200;
			16'h2ffe: y = 16'h200;
			16'h2fff: y = 16'h200;
			16'h3000: y = 16'h200;
			16'h3001: y = 16'h200;
			16'h3002: y = 16'h200;
			16'h3003: y = 16'h200;
			16'h3004: y = 16'h200;
			16'h3005: y = 16'h200;
			16'h3006: y = 16'h200;
			16'h3007: y = 16'h200;
			16'h3008: y = 16'h200;
			16'h3009: y = 16'h200;
			16'h300a: y = 16'h200;
			16'h300b: y = 16'h200;
			16'h300c: y = 16'h200;
			16'h300d: y = 16'h200;
			16'h300e: y = 16'h200;
			16'h300f: y = 16'h200;
			16'h3010: y = 16'h200;
			16'h3011: y = 16'h200;
			16'h3012: y = 16'h200;
			16'h3013: y = 16'h200;
			16'h3014: y = 16'h200;
			16'h3015: y = 16'h200;
			16'h3016: y = 16'h200;
			16'h3017: y = 16'h200;
			16'h3018: y = 16'h200;
			16'h3019: y = 16'h200;
			16'h301a: y = 16'h200;
			16'h301b: y = 16'h200;
			16'h301c: y = 16'h200;
			16'h301d: y = 16'h200;
			16'h301e: y = 16'h200;
			16'h301f: y = 16'h200;
			16'h3020: y = 16'h200;
			16'h3021: y = 16'h200;
			16'h3022: y = 16'h200;
			16'h3023: y = 16'h200;
			16'h3024: y = 16'h200;
			16'h3025: y = 16'h200;
			16'h3026: y = 16'h200;
			16'h3027: y = 16'h200;
			16'h3028: y = 16'h200;
			16'h3029: y = 16'h200;
			16'h302a: y = 16'h200;
			16'h302b: y = 16'h200;
			16'h302c: y = 16'h200;
			16'h302d: y = 16'h200;
			16'h302e: y = 16'h200;
			16'h302f: y = 16'h200;
			16'h3030: y = 16'h200;
			16'h3031: y = 16'h200;
			16'h3032: y = 16'h200;
			16'h3033: y = 16'h200;
			16'h3034: y = 16'h200;
			16'h3035: y = 16'h200;
			16'h3036: y = 16'h200;
			16'h3037: y = 16'h200;
			16'h3038: y = 16'h200;
			16'h3039: y = 16'h200;
			16'h303a: y = 16'h200;
			16'h303b: y = 16'h200;
			16'h303c: y = 16'h200;
			16'h303d: y = 16'h200;
			16'h303e: y = 16'h200;
			16'h303f: y = 16'h200;
			16'h3040: y = 16'h200;
			16'h3041: y = 16'h200;
			16'h3042: y = 16'h200;
			16'h3043: y = 16'h200;
			16'h3044: y = 16'h200;
			16'h3045: y = 16'h200;
			16'h3046: y = 16'h200;
			16'h3047: y = 16'h200;
			16'h3048: y = 16'h200;
			16'h3049: y = 16'h200;
			16'h304a: y = 16'h200;
			16'h304b: y = 16'h200;
			16'h304c: y = 16'h200;
			16'h304d: y = 16'h200;
			16'h304e: y = 16'h200;
			16'h304f: y = 16'h200;
			16'h3050: y = 16'h200;
			16'h3051: y = 16'h200;
			16'h3052: y = 16'h200;
			16'h3053: y = 16'h200;
			16'h3054: y = 16'h200;
			16'h3055: y = 16'h200;
			16'h3056: y = 16'h200;
			16'h3057: y = 16'h200;
			16'h3058: y = 16'h200;
			16'h3059: y = 16'h200;
			16'h305a: y = 16'h200;
			16'h305b: y = 16'h200;
			16'h305c: y = 16'h200;
			16'h305d: y = 16'h200;
			16'h305e: y = 16'h200;
			16'h305f: y = 16'h200;
			16'h3060: y = 16'h200;
			16'h3061: y = 16'h200;
			16'h3062: y = 16'h200;
			16'h3063: y = 16'h200;
			16'h3064: y = 16'h200;
			16'h3065: y = 16'h200;
			16'h3066: y = 16'h200;
			16'h3067: y = 16'h200;
			16'h3068: y = 16'h200;
			16'h3069: y = 16'h200;
			16'h306a: y = 16'h200;
			16'h306b: y = 16'h200;
			16'h306c: y = 16'h200;
			16'h306d: y = 16'h200;
			16'h306e: y = 16'h200;
			16'h306f: y = 16'h200;
			16'h3070: y = 16'h200;
			16'h3071: y = 16'h200;
			16'h3072: y = 16'h200;
			16'h3073: y = 16'h200;
			16'h3074: y = 16'h200;
			16'h3075: y = 16'h200;
			16'h3076: y = 16'h200;
			16'h3077: y = 16'h200;
			16'h3078: y = 16'h200;
			16'h3079: y = 16'h200;
			16'h307a: y = 16'h200;
			16'h307b: y = 16'h200;
			16'h307c: y = 16'h200;
			16'h307d: y = 16'h200;
			16'h307e: y = 16'h200;
			16'h307f: y = 16'h200;
			16'h3080: y = 16'h200;
			16'h3081: y = 16'h200;
			16'h3082: y = 16'h200;
			16'h3083: y = 16'h200;
			16'h3084: y = 16'h200;
			16'h3085: y = 16'h200;
			16'h3086: y = 16'h200;
			16'h3087: y = 16'h200;
			16'h3088: y = 16'h200;
			16'h3089: y = 16'h200;
			16'h308a: y = 16'h200;
			16'h308b: y = 16'h200;
			16'h308c: y = 16'h200;
			16'h308d: y = 16'h200;
			16'h308e: y = 16'h200;
			16'h308f: y = 16'h200;
			16'h3090: y = 16'h200;
			16'h3091: y = 16'h200;
			16'h3092: y = 16'h200;
			16'h3093: y = 16'h200;
			16'h3094: y = 16'h200;
			16'h3095: y = 16'h200;
			16'h3096: y = 16'h200;
			16'h3097: y = 16'h200;
			16'h3098: y = 16'h200;
			16'h3099: y = 16'h200;
			16'h309a: y = 16'h200;
			16'h309b: y = 16'h200;
			16'h309c: y = 16'h200;
			16'h309d: y = 16'h200;
			16'h309e: y = 16'h200;
			16'h309f: y = 16'h200;
			16'h30a0: y = 16'h200;
			16'h30a1: y = 16'h200;
			16'h30a2: y = 16'h200;
			16'h30a3: y = 16'h200;
			16'h30a4: y = 16'h200;
			16'h30a5: y = 16'h200;
			16'h30a6: y = 16'h200;
			16'h30a7: y = 16'h200;
			16'h30a8: y = 16'h200;
			16'h30a9: y = 16'h200;
			16'h30aa: y = 16'h200;
			16'h30ab: y = 16'h200;
			16'h30ac: y = 16'h200;
			16'h30ad: y = 16'h200;
			16'h30ae: y = 16'h200;
			16'h30af: y = 16'h200;
			16'h30b0: y = 16'h200;
			16'h30b1: y = 16'h200;
			16'h30b2: y = 16'h200;
			16'h30b3: y = 16'h200;
			16'h30b4: y = 16'h200;
			16'h30b5: y = 16'h200;
			16'h30b6: y = 16'h200;
			16'h30b7: y = 16'h200;
			16'h30b8: y = 16'h200;
			16'h30b9: y = 16'h200;
			16'h30ba: y = 16'h200;
			16'h30bb: y = 16'h200;
			16'h30bc: y = 16'h200;
			16'h30bd: y = 16'h200;
			16'h30be: y = 16'h200;
			16'h30bf: y = 16'h200;
			16'h30c0: y = 16'h200;
			16'h30c1: y = 16'h200;
			16'h30c2: y = 16'h200;
			16'h30c3: y = 16'h200;
			16'h30c4: y = 16'h200;
			16'h30c5: y = 16'h200;
			16'h30c6: y = 16'h200;
			16'h30c7: y = 16'h200;
			16'h30c8: y = 16'h200;
			16'h30c9: y = 16'h200;
			16'h30ca: y = 16'h200;
			16'h30cb: y = 16'h200;
			16'h30cc: y = 16'h200;
			16'h30cd: y = 16'h200;
			16'h30ce: y = 16'h200;
			16'h30cf: y = 16'h200;
			16'h30d0: y = 16'h200;
			16'h30d1: y = 16'h200;
			16'h30d2: y = 16'h200;
			16'h30d3: y = 16'h200;
			16'h30d4: y = 16'h200;
			16'h30d5: y = 16'h200;
			16'h30d6: y = 16'h200;
			16'h30d7: y = 16'h200;
			16'h30d8: y = 16'h200;
			16'h30d9: y = 16'h200;
			16'h30da: y = 16'h200;
			16'h30db: y = 16'h200;
			16'h30dc: y = 16'h200;
			16'h30dd: y = 16'h200;
			16'h30de: y = 16'h200;
			16'h30df: y = 16'h200;
			16'h30e0: y = 16'h200;
			16'h30e1: y = 16'h200;
			16'h30e2: y = 16'h200;
			16'h30e3: y = 16'h200;
			16'h30e4: y = 16'h200;
			16'h30e5: y = 16'h200;
			16'h30e6: y = 16'h200;
			16'h30e7: y = 16'h200;
			16'h30e8: y = 16'h200;
			16'h30e9: y = 16'h200;
			16'h30ea: y = 16'h200;
			16'h30eb: y = 16'h200;
			16'h30ec: y = 16'h200;
			16'h30ed: y = 16'h200;
			16'h30ee: y = 16'h200;
			16'h30ef: y = 16'h200;
			16'h30f0: y = 16'h200;
			16'h30f1: y = 16'h200;
			16'h30f2: y = 16'h200;
			16'h30f3: y = 16'h200;
			16'h30f4: y = 16'h200;
			16'h30f5: y = 16'h200;
			16'h30f6: y = 16'h200;
			16'h30f7: y = 16'h200;
			16'h30f8: y = 16'h200;
			16'h30f9: y = 16'h200;
			16'h30fa: y = 16'h200;
			16'h30fb: y = 16'h200;
			16'h30fc: y = 16'h200;
			16'h30fd: y = 16'h200;
			16'h30fe: y = 16'h200;
			16'h30ff: y = 16'h200;
			16'h3100: y = 16'h200;
			16'h3101: y = 16'h200;
			16'h3102: y = 16'h200;
			16'h3103: y = 16'h200;
			16'h3104: y = 16'h200;
			16'h3105: y = 16'h200;
			16'h3106: y = 16'h200;
			16'h3107: y = 16'h200;
			16'h3108: y = 16'h200;
			16'h3109: y = 16'h200;
			16'h310a: y = 16'h200;
			16'h310b: y = 16'h200;
			16'h310c: y = 16'h200;
			16'h310d: y = 16'h200;
			16'h310e: y = 16'h200;
			16'h310f: y = 16'h200;
			16'h3110: y = 16'h200;
			16'h3111: y = 16'h200;
			16'h3112: y = 16'h200;
			16'h3113: y = 16'h200;
			16'h3114: y = 16'h200;
			16'h3115: y = 16'h200;
			16'h3116: y = 16'h200;
			16'h3117: y = 16'h200;
			16'h3118: y = 16'h200;
			16'h3119: y = 16'h200;
			16'h311a: y = 16'h200;
			16'h311b: y = 16'h200;
			16'h311c: y = 16'h200;
			16'h311d: y = 16'h200;
			16'h311e: y = 16'h200;
			16'h311f: y = 16'h200;
			16'h3120: y = 16'h200;
			16'h3121: y = 16'h200;
			16'h3122: y = 16'h200;
			16'h3123: y = 16'h200;
			16'h3124: y = 16'h200;
			16'h3125: y = 16'h200;
			16'h3126: y = 16'h200;
			16'h3127: y = 16'h200;
			16'h3128: y = 16'h200;
			16'h3129: y = 16'h200;
			16'h312a: y = 16'h200;
			16'h312b: y = 16'h200;
			16'h312c: y = 16'h200;
			16'h312d: y = 16'h200;
			16'h312e: y = 16'h200;
			16'h312f: y = 16'h200;
			16'h3130: y = 16'h200;
			16'h3131: y = 16'h200;
			16'h3132: y = 16'h200;
			16'h3133: y = 16'h200;
			16'h3134: y = 16'h200;
			16'h3135: y = 16'h200;
			16'h3136: y = 16'h200;
			16'h3137: y = 16'h200;
			16'h3138: y = 16'h200;
			16'h3139: y = 16'h200;
			16'h313a: y = 16'h200;
			16'h313b: y = 16'h200;
			16'h313c: y = 16'h200;
			16'h313d: y = 16'h200;
			16'h313e: y = 16'h200;
			16'h313f: y = 16'h200;
			16'h3140: y = 16'h200;
			16'h3141: y = 16'h200;
			16'h3142: y = 16'h200;
			16'h3143: y = 16'h200;
			16'h3144: y = 16'h200;
			16'h3145: y = 16'h200;
			16'h3146: y = 16'h200;
			16'h3147: y = 16'h200;
			16'h3148: y = 16'h200;
			16'h3149: y = 16'h200;
			16'h314a: y = 16'h200;
			16'h314b: y = 16'h200;
			16'h314c: y = 16'h200;
			16'h314d: y = 16'h200;
			16'h314e: y = 16'h200;
			16'h314f: y = 16'h200;
			16'h3150: y = 16'h200;
			16'h3151: y = 16'h200;
			16'h3152: y = 16'h200;
			16'h3153: y = 16'h200;
			16'h3154: y = 16'h200;
			16'h3155: y = 16'h200;
			16'h3156: y = 16'h200;
			16'h3157: y = 16'h200;
			16'h3158: y = 16'h200;
			16'h3159: y = 16'h200;
			16'h315a: y = 16'h200;
			16'h315b: y = 16'h200;
			16'h315c: y = 16'h200;
			16'h315d: y = 16'h200;
			16'h315e: y = 16'h200;
			16'h315f: y = 16'h200;
			16'h3160: y = 16'h200;
			16'h3161: y = 16'h200;
			16'h3162: y = 16'h200;
			16'h3163: y = 16'h200;
			16'h3164: y = 16'h200;
			16'h3165: y = 16'h200;
			16'h3166: y = 16'h200;
			16'h3167: y = 16'h200;
			16'h3168: y = 16'h200;
			16'h3169: y = 16'h200;
			16'h316a: y = 16'h200;
			16'h316b: y = 16'h200;
			16'h316c: y = 16'h200;
			16'h316d: y = 16'h200;
			16'h316e: y = 16'h200;
			16'h316f: y = 16'h200;
			16'h3170: y = 16'h200;
			16'h3171: y = 16'h200;
			16'h3172: y = 16'h200;
			16'h3173: y = 16'h200;
			16'h3174: y = 16'h200;
			16'h3175: y = 16'h200;
			16'h3176: y = 16'h200;
			16'h3177: y = 16'h200;
			16'h3178: y = 16'h200;
			16'h3179: y = 16'h200;
			16'h317a: y = 16'h200;
			16'h317b: y = 16'h200;
			16'h317c: y = 16'h200;
			16'h317d: y = 16'h200;
			16'h317e: y = 16'h200;
			16'h317f: y = 16'h200;
			16'h3180: y = 16'h200;
			16'h3181: y = 16'h200;
			16'h3182: y = 16'h200;
			16'h3183: y = 16'h200;
			16'h3184: y = 16'h200;
			16'h3185: y = 16'h200;
			16'h3186: y = 16'h200;
			16'h3187: y = 16'h200;
			16'h3188: y = 16'h200;
			16'h3189: y = 16'h200;
			16'h318a: y = 16'h200;
			16'h318b: y = 16'h200;
			16'h318c: y = 16'h200;
			16'h318d: y = 16'h200;
			16'h318e: y = 16'h200;
			16'h318f: y = 16'h200;
			16'h3190: y = 16'h200;
			16'h3191: y = 16'h200;
			16'h3192: y = 16'h200;
			16'h3193: y = 16'h200;
			16'h3194: y = 16'h200;
			16'h3195: y = 16'h200;
			16'h3196: y = 16'h200;
			16'h3197: y = 16'h200;
			16'h3198: y = 16'h200;
			16'h3199: y = 16'h200;
			16'h319a: y = 16'h200;
			16'h319b: y = 16'h200;
			16'h319c: y = 16'h200;
			16'h319d: y = 16'h200;
			16'h319e: y = 16'h200;
			16'h319f: y = 16'h200;
			16'h31a0: y = 16'h200;
			16'h31a1: y = 16'h200;
			16'h31a2: y = 16'h200;
			16'h31a3: y = 16'h200;
			16'h31a4: y = 16'h200;
			16'h31a5: y = 16'h200;
			16'h31a6: y = 16'h200;
			16'h31a7: y = 16'h200;
			16'h31a8: y = 16'h200;
			16'h31a9: y = 16'h200;
			16'h31aa: y = 16'h200;
			16'h31ab: y = 16'h200;
			16'h31ac: y = 16'h200;
			16'h31ad: y = 16'h200;
			16'h31ae: y = 16'h200;
			16'h31af: y = 16'h200;
			16'h31b0: y = 16'h200;
			16'h31b1: y = 16'h200;
			16'h31b2: y = 16'h200;
			16'h31b3: y = 16'h200;
			16'h31b4: y = 16'h200;
			16'h31b5: y = 16'h200;
			16'h31b6: y = 16'h200;
			16'h31b7: y = 16'h200;
			16'h31b8: y = 16'h200;
			16'h31b9: y = 16'h200;
			16'h31ba: y = 16'h200;
			16'h31bb: y = 16'h200;
			16'h31bc: y = 16'h200;
			16'h31bd: y = 16'h200;
			16'h31be: y = 16'h200;
			16'h31bf: y = 16'h200;
			16'h31c0: y = 16'h200;
			16'h31c1: y = 16'h200;
			16'h31c2: y = 16'h200;
			16'h31c3: y = 16'h200;
			16'h31c4: y = 16'h200;
			16'h31c5: y = 16'h200;
			16'h31c6: y = 16'h200;
			16'h31c7: y = 16'h200;
			16'h31c8: y = 16'h200;
			16'h31c9: y = 16'h200;
			16'h31ca: y = 16'h200;
			16'h31cb: y = 16'h200;
			16'h31cc: y = 16'h200;
			16'h31cd: y = 16'h200;
			16'h31ce: y = 16'h200;
			16'h31cf: y = 16'h200;
			16'h31d0: y = 16'h200;
			16'h31d1: y = 16'h200;
			16'h31d2: y = 16'h200;
			16'h31d3: y = 16'h200;
			16'h31d4: y = 16'h200;
			16'h31d5: y = 16'h200;
			16'h31d6: y = 16'h200;
			16'h31d7: y = 16'h200;
			16'h31d8: y = 16'h200;
			16'h31d9: y = 16'h200;
			16'h31da: y = 16'h200;
			16'h31db: y = 16'h200;
			16'h31dc: y = 16'h200;
			16'h31dd: y = 16'h200;
			16'h31de: y = 16'h200;
			16'h31df: y = 16'h200;
			16'h31e0: y = 16'h200;
			16'h31e1: y = 16'h200;
			16'h31e2: y = 16'h200;
			16'h31e3: y = 16'h200;
			16'h31e4: y = 16'h200;
			16'h31e5: y = 16'h200;
			16'h31e6: y = 16'h200;
			16'h31e7: y = 16'h200;
			16'h31e8: y = 16'h200;
			16'h31e9: y = 16'h200;
			16'h31ea: y = 16'h200;
			16'h31eb: y = 16'h200;
			16'h31ec: y = 16'h200;
			16'h31ed: y = 16'h200;
			16'h31ee: y = 16'h200;
			16'h31ef: y = 16'h200;
			16'h31f0: y = 16'h200;
			16'h31f1: y = 16'h200;
			16'h31f2: y = 16'h200;
			16'h31f3: y = 16'h200;
			16'h31f4: y = 16'h200;
			16'h31f5: y = 16'h200;
			16'h31f6: y = 16'h200;
			16'h31f7: y = 16'h200;
			16'h31f8: y = 16'h200;
			16'h31f9: y = 16'h200;
			16'h31fa: y = 16'h200;
			16'h31fb: y = 16'h200;
			16'h31fc: y = 16'h200;
			16'h31fd: y = 16'h200;
			16'h31fe: y = 16'h200;
			16'h31ff: y = 16'h200;
			16'h3200: y = 16'h200;
			16'h3201: y = 16'h200;
			16'h3202: y = 16'h200;
			16'h3203: y = 16'h200;
			16'h3204: y = 16'h200;
			16'h3205: y = 16'h200;
			16'h3206: y = 16'h200;
			16'h3207: y = 16'h200;
			16'h3208: y = 16'h200;
			16'h3209: y = 16'h200;
			16'h320a: y = 16'h200;
			16'h320b: y = 16'h200;
			16'h320c: y = 16'h200;
			16'h320d: y = 16'h200;
			16'h320e: y = 16'h200;
			16'h320f: y = 16'h200;
			16'h3210: y = 16'h200;
			16'h3211: y = 16'h200;
			16'h3212: y = 16'h200;
			16'h3213: y = 16'h200;
			16'h3214: y = 16'h200;
			16'h3215: y = 16'h200;
			16'h3216: y = 16'h200;
			16'h3217: y = 16'h200;
			16'h3218: y = 16'h200;
			16'h3219: y = 16'h200;
			16'h321a: y = 16'h200;
			16'h321b: y = 16'h200;
			16'h321c: y = 16'h200;
			16'h321d: y = 16'h200;
			16'h321e: y = 16'h200;
			16'h321f: y = 16'h200;
			16'h3220: y = 16'h200;
			16'h3221: y = 16'h200;
			16'h3222: y = 16'h200;
			16'h3223: y = 16'h200;
			16'h3224: y = 16'h200;
			16'h3225: y = 16'h200;
			16'h3226: y = 16'h200;
			16'h3227: y = 16'h200;
			16'h3228: y = 16'h200;
			16'h3229: y = 16'h200;
			16'h322a: y = 16'h200;
			16'h322b: y = 16'h200;
			16'h322c: y = 16'h200;
			16'h322d: y = 16'h200;
			16'h322e: y = 16'h200;
			16'h322f: y = 16'h200;
			16'h3230: y = 16'h200;
			16'h3231: y = 16'h200;
			16'h3232: y = 16'h200;
			16'h3233: y = 16'h200;
			16'h3234: y = 16'h200;
			16'h3235: y = 16'h200;
			16'h3236: y = 16'h200;
			16'h3237: y = 16'h200;
			16'h3238: y = 16'h200;
			16'h3239: y = 16'h200;
			16'h323a: y = 16'h200;
			16'h323b: y = 16'h200;
			16'h323c: y = 16'h200;
			16'h323d: y = 16'h200;
			16'h323e: y = 16'h200;
			16'h323f: y = 16'h200;
			16'h3240: y = 16'h200;
			16'h3241: y = 16'h200;
			16'h3242: y = 16'h200;
			16'h3243: y = 16'h200;
			16'h3244: y = 16'h200;
			16'h3245: y = 16'h200;
			16'h3246: y = 16'h200;
			16'h3247: y = 16'h200;
			16'h3248: y = 16'h200;
			16'h3249: y = 16'h200;
			16'h324a: y = 16'h200;
			16'h324b: y = 16'h200;
			16'h324c: y = 16'h200;
			16'h324d: y = 16'h200;
			16'h324e: y = 16'h200;
			16'h324f: y = 16'h200;
			16'h3250: y = 16'h200;
			16'h3251: y = 16'h200;
			16'h3252: y = 16'h200;
			16'h3253: y = 16'h200;
			16'h3254: y = 16'h200;
			16'h3255: y = 16'h200;
			16'h3256: y = 16'h200;
			16'h3257: y = 16'h200;
			16'h3258: y = 16'h200;
			16'h3259: y = 16'h200;
			16'h325a: y = 16'h200;
			16'h325b: y = 16'h200;
			16'h325c: y = 16'h200;
			16'h325d: y = 16'h200;
			16'h325e: y = 16'h200;
			16'h325f: y = 16'h200;
			16'h3260: y = 16'h200;
			16'h3261: y = 16'h200;
			16'h3262: y = 16'h200;
			16'h3263: y = 16'h200;
			16'h3264: y = 16'h200;
			16'h3265: y = 16'h200;
			16'h3266: y = 16'h200;
			16'h3267: y = 16'h200;
			16'h3268: y = 16'h200;
			16'h3269: y = 16'h200;
			16'h326a: y = 16'h200;
			16'h326b: y = 16'h200;
			16'h326c: y = 16'h200;
			16'h326d: y = 16'h200;
			16'h326e: y = 16'h200;
			16'h326f: y = 16'h200;
			16'h3270: y = 16'h200;
			16'h3271: y = 16'h200;
			16'h3272: y = 16'h200;
			16'h3273: y = 16'h200;
			16'h3274: y = 16'h200;
			16'h3275: y = 16'h200;
			16'h3276: y = 16'h200;
			16'h3277: y = 16'h200;
			16'h3278: y = 16'h200;
			16'h3279: y = 16'h200;
			16'h327a: y = 16'h200;
			16'h327b: y = 16'h200;
			16'h327c: y = 16'h200;
			16'h327d: y = 16'h200;
			16'h327e: y = 16'h200;
			16'h327f: y = 16'h200;
			16'h3280: y = 16'h200;
			16'h3281: y = 16'h200;
			16'h3282: y = 16'h200;
			16'h3283: y = 16'h200;
			16'h3284: y = 16'h200;
			16'h3285: y = 16'h200;
			16'h3286: y = 16'h200;
			16'h3287: y = 16'h200;
			16'h3288: y = 16'h200;
			16'h3289: y = 16'h200;
			16'h328a: y = 16'h200;
			16'h328b: y = 16'h200;
			16'h328c: y = 16'h200;
			16'h328d: y = 16'h200;
			16'h328e: y = 16'h200;
			16'h328f: y = 16'h200;
			16'h3290: y = 16'h200;
			16'h3291: y = 16'h200;
			16'h3292: y = 16'h200;
			16'h3293: y = 16'h200;
			16'h3294: y = 16'h200;
			16'h3295: y = 16'h200;
			16'h3296: y = 16'h200;
			16'h3297: y = 16'h200;
			16'h3298: y = 16'h200;
			16'h3299: y = 16'h200;
			16'h329a: y = 16'h200;
			16'h329b: y = 16'h200;
			16'h329c: y = 16'h200;
			16'h329d: y = 16'h200;
			16'h329e: y = 16'h200;
			16'h329f: y = 16'h200;
			16'h32a0: y = 16'h200;
			16'h32a1: y = 16'h200;
			16'h32a2: y = 16'h200;
			16'h32a3: y = 16'h200;
			16'h32a4: y = 16'h200;
			16'h32a5: y = 16'h200;
			16'h32a6: y = 16'h200;
			16'h32a7: y = 16'h200;
			16'h32a8: y = 16'h200;
			16'h32a9: y = 16'h200;
			16'h32aa: y = 16'h200;
			16'h32ab: y = 16'h200;
			16'h32ac: y = 16'h200;
			16'h32ad: y = 16'h200;
			16'h32ae: y = 16'h200;
			16'h32af: y = 16'h200;
			16'h32b0: y = 16'h200;
			16'h32b1: y = 16'h200;
			16'h32b2: y = 16'h200;
			16'h32b3: y = 16'h200;
			16'h32b4: y = 16'h200;
			16'h32b5: y = 16'h200;
			16'h32b6: y = 16'h200;
			16'h32b7: y = 16'h200;
			16'h32b8: y = 16'h200;
			16'h32b9: y = 16'h200;
			16'h32ba: y = 16'h200;
			16'h32bb: y = 16'h200;
			16'h32bc: y = 16'h200;
			16'h32bd: y = 16'h200;
			16'h32be: y = 16'h200;
			16'h32bf: y = 16'h200;
			16'h32c0: y = 16'h200;
			16'h32c1: y = 16'h200;
			16'h32c2: y = 16'h200;
			16'h32c3: y = 16'h200;
			16'h32c4: y = 16'h200;
			16'h32c5: y = 16'h200;
			16'h32c6: y = 16'h200;
			16'h32c7: y = 16'h200;
			16'h32c8: y = 16'h200;
			16'h32c9: y = 16'h200;
			16'h32ca: y = 16'h200;
			16'h32cb: y = 16'h200;
			16'h32cc: y = 16'h200;
			16'h32cd: y = 16'h200;
			16'h32ce: y = 16'h200;
			16'h32cf: y = 16'h200;
			16'h32d0: y = 16'h200;
			16'h32d1: y = 16'h200;
			16'h32d2: y = 16'h200;
			16'h32d3: y = 16'h200;
			16'h32d4: y = 16'h200;
			16'h32d5: y = 16'h200;
			16'h32d6: y = 16'h200;
			16'h32d7: y = 16'h200;
			16'h32d8: y = 16'h200;
			16'h32d9: y = 16'h200;
			16'h32da: y = 16'h200;
			16'h32db: y = 16'h200;
			16'h32dc: y = 16'h200;
			16'h32dd: y = 16'h200;
			16'h32de: y = 16'h200;
			16'h32df: y = 16'h200;
			16'h32e0: y = 16'h200;
			16'h32e1: y = 16'h200;
			16'h32e2: y = 16'h200;
			16'h32e3: y = 16'h200;
			16'h32e4: y = 16'h200;
			16'h32e5: y = 16'h200;
			16'h32e6: y = 16'h200;
			16'h32e7: y = 16'h200;
			16'h32e8: y = 16'h200;
			16'h32e9: y = 16'h200;
			16'h32ea: y = 16'h200;
			16'h32eb: y = 16'h200;
			16'h32ec: y = 16'h200;
			16'h32ed: y = 16'h200;
			16'h32ee: y = 16'h200;
			16'h32ef: y = 16'h200;
			16'h32f0: y = 16'h200;
			16'h32f1: y = 16'h200;
			16'h32f2: y = 16'h200;
			16'h32f3: y = 16'h200;
			16'h32f4: y = 16'h200;
			16'h32f5: y = 16'h200;
			16'h32f6: y = 16'h200;
			16'h32f7: y = 16'h200;
			16'h32f8: y = 16'h200;
			16'h32f9: y = 16'h200;
			16'h32fa: y = 16'h200;
			16'h32fb: y = 16'h200;
			16'h32fc: y = 16'h200;
			16'h32fd: y = 16'h200;
			16'h32fe: y = 16'h200;
			16'h32ff: y = 16'h200;
			16'h3300: y = 16'h200;
			16'h3301: y = 16'h200;
			16'h3302: y = 16'h200;
			16'h3303: y = 16'h200;
			16'h3304: y = 16'h200;
			16'h3305: y = 16'h200;
			16'h3306: y = 16'h200;
			16'h3307: y = 16'h200;
			16'h3308: y = 16'h200;
			16'h3309: y = 16'h200;
			16'h330a: y = 16'h200;
			16'h330b: y = 16'h200;
			16'h330c: y = 16'h200;
			16'h330d: y = 16'h200;
			16'h330e: y = 16'h200;
			16'h330f: y = 16'h200;
			16'h3310: y = 16'h200;
			16'h3311: y = 16'h200;
			16'h3312: y = 16'h200;
			16'h3313: y = 16'h200;
			16'h3314: y = 16'h200;
			16'h3315: y = 16'h200;
			16'h3316: y = 16'h200;
			16'h3317: y = 16'h200;
			16'h3318: y = 16'h200;
			16'h3319: y = 16'h200;
			16'h331a: y = 16'h200;
			16'h331b: y = 16'h200;
			16'h331c: y = 16'h200;
			16'h331d: y = 16'h200;
			16'h331e: y = 16'h200;
			16'h331f: y = 16'h200;
			16'h3320: y = 16'h200;
			16'h3321: y = 16'h200;
			16'h3322: y = 16'h200;
			16'h3323: y = 16'h200;
			16'h3324: y = 16'h200;
			16'h3325: y = 16'h200;
			16'h3326: y = 16'h200;
			16'h3327: y = 16'h200;
			16'h3328: y = 16'h200;
			16'h3329: y = 16'h200;
			16'h332a: y = 16'h200;
			16'h332b: y = 16'h200;
			16'h332c: y = 16'h200;
			16'h332d: y = 16'h200;
			16'h332e: y = 16'h200;
			16'h332f: y = 16'h200;
			16'h3330: y = 16'h200;
			16'h3331: y = 16'h200;
			16'h3332: y = 16'h200;
			16'h3333: y = 16'h200;
			16'h3334: y = 16'h200;
			16'h3335: y = 16'h200;
			16'h3336: y = 16'h200;
			16'h3337: y = 16'h200;
			16'h3338: y = 16'h200;
			16'h3339: y = 16'h200;
			16'h333a: y = 16'h200;
			16'h333b: y = 16'h200;
			16'h333c: y = 16'h200;
			16'h333d: y = 16'h200;
			16'h333e: y = 16'h200;
			16'h333f: y = 16'h200;
			16'h3340: y = 16'h200;
			16'h3341: y = 16'h200;
			16'h3342: y = 16'h200;
			16'h3343: y = 16'h200;
			16'h3344: y = 16'h200;
			16'h3345: y = 16'h200;
			16'h3346: y = 16'h200;
			16'h3347: y = 16'h200;
			16'h3348: y = 16'h200;
			16'h3349: y = 16'h200;
			16'h334a: y = 16'h200;
			16'h334b: y = 16'h200;
			16'h334c: y = 16'h200;
			16'h334d: y = 16'h200;
			16'h334e: y = 16'h200;
			16'h334f: y = 16'h200;
			16'h3350: y = 16'h200;
			16'h3351: y = 16'h200;
			16'h3352: y = 16'h200;
			16'h3353: y = 16'h200;
			16'h3354: y = 16'h200;
			16'h3355: y = 16'h200;
			16'h3356: y = 16'h200;
			16'h3357: y = 16'h200;
			16'h3358: y = 16'h200;
			16'h3359: y = 16'h200;
			16'h335a: y = 16'h200;
			16'h335b: y = 16'h200;
			16'h335c: y = 16'h200;
			16'h335d: y = 16'h200;
			16'h335e: y = 16'h200;
			16'h335f: y = 16'h200;
			16'h3360: y = 16'h200;
			16'h3361: y = 16'h200;
			16'h3362: y = 16'h200;
			16'h3363: y = 16'h200;
			16'h3364: y = 16'h200;
			16'h3365: y = 16'h200;
			16'h3366: y = 16'h200;
			16'h3367: y = 16'h200;
			16'h3368: y = 16'h200;
			16'h3369: y = 16'h200;
			16'h336a: y = 16'h200;
			16'h336b: y = 16'h200;
			16'h336c: y = 16'h200;
			16'h336d: y = 16'h200;
			16'h336e: y = 16'h200;
			16'h336f: y = 16'h200;
			16'h3370: y = 16'h200;
			16'h3371: y = 16'h200;
			16'h3372: y = 16'h200;
			16'h3373: y = 16'h200;
			16'h3374: y = 16'h200;
			16'h3375: y = 16'h200;
			16'h3376: y = 16'h200;
			16'h3377: y = 16'h200;
			16'h3378: y = 16'h200;
			16'h3379: y = 16'h200;
			16'h337a: y = 16'h200;
			16'h337b: y = 16'h200;
			16'h337c: y = 16'h200;
			16'h337d: y = 16'h200;
			16'h337e: y = 16'h200;
			16'h337f: y = 16'h200;
			16'h3380: y = 16'h200;
			16'h3381: y = 16'h200;
			16'h3382: y = 16'h200;
			16'h3383: y = 16'h200;
			16'h3384: y = 16'h200;
			16'h3385: y = 16'h200;
			16'h3386: y = 16'h200;
			16'h3387: y = 16'h200;
			16'h3388: y = 16'h200;
			16'h3389: y = 16'h200;
			16'h338a: y = 16'h200;
			16'h338b: y = 16'h200;
			16'h338c: y = 16'h200;
			16'h338d: y = 16'h200;
			16'h338e: y = 16'h200;
			16'h338f: y = 16'h200;
			16'h3390: y = 16'h200;
			16'h3391: y = 16'h200;
			16'h3392: y = 16'h200;
			16'h3393: y = 16'h200;
			16'h3394: y = 16'h200;
			16'h3395: y = 16'h200;
			16'h3396: y = 16'h200;
			16'h3397: y = 16'h200;
			16'h3398: y = 16'h200;
			16'h3399: y = 16'h200;
			16'h339a: y = 16'h200;
			16'h339b: y = 16'h200;
			16'h339c: y = 16'h200;
			16'h339d: y = 16'h200;
			16'h339e: y = 16'h200;
			16'h339f: y = 16'h200;
			16'h33a0: y = 16'h200;
			16'h33a1: y = 16'h200;
			16'h33a2: y = 16'h200;
			16'h33a3: y = 16'h200;
			16'h33a4: y = 16'h200;
			16'h33a5: y = 16'h200;
			16'h33a6: y = 16'h200;
			16'h33a7: y = 16'h200;
			16'h33a8: y = 16'h200;
			16'h33a9: y = 16'h200;
			16'h33aa: y = 16'h200;
			16'h33ab: y = 16'h200;
			16'h33ac: y = 16'h200;
			16'h33ad: y = 16'h200;
			16'h33ae: y = 16'h200;
			16'h33af: y = 16'h200;
			16'h33b0: y = 16'h200;
			16'h33b1: y = 16'h200;
			16'h33b2: y = 16'h200;
			16'h33b3: y = 16'h200;
			16'h33b4: y = 16'h200;
			16'h33b5: y = 16'h200;
			16'h33b6: y = 16'h200;
			16'h33b7: y = 16'h200;
			16'h33b8: y = 16'h200;
			16'h33b9: y = 16'h200;
			16'h33ba: y = 16'h200;
			16'h33bb: y = 16'h200;
			16'h33bc: y = 16'h200;
			16'h33bd: y = 16'h200;
			16'h33be: y = 16'h200;
			16'h33bf: y = 16'h200;
			16'h33c0: y = 16'h200;
			16'h33c1: y = 16'h200;
			16'h33c2: y = 16'h200;
			16'h33c3: y = 16'h200;
			16'h33c4: y = 16'h200;
			16'h33c5: y = 16'h200;
			16'h33c6: y = 16'h200;
			16'h33c7: y = 16'h200;
			16'h33c8: y = 16'h200;
			16'h33c9: y = 16'h200;
			16'h33ca: y = 16'h200;
			16'h33cb: y = 16'h200;
			16'h33cc: y = 16'h200;
			16'h33cd: y = 16'h200;
			16'h33ce: y = 16'h200;
			16'h33cf: y = 16'h200;
			16'h33d0: y = 16'h200;
			16'h33d1: y = 16'h200;
			16'h33d2: y = 16'h200;
			16'h33d3: y = 16'h200;
			16'h33d4: y = 16'h200;
			16'h33d5: y = 16'h200;
			16'h33d6: y = 16'h200;
			16'h33d7: y = 16'h200;
			16'h33d8: y = 16'h200;
			16'h33d9: y = 16'h200;
			16'h33da: y = 16'h200;
			16'h33db: y = 16'h200;
			16'h33dc: y = 16'h200;
			16'h33dd: y = 16'h200;
			16'h33de: y = 16'h200;
			16'h33df: y = 16'h200;
			16'h33e0: y = 16'h200;
			16'h33e1: y = 16'h200;
			16'h33e2: y = 16'h200;
			16'h33e3: y = 16'h200;
			16'h33e4: y = 16'h200;
			16'h33e5: y = 16'h200;
			16'h33e6: y = 16'h200;
			16'h33e7: y = 16'h200;
			16'h33e8: y = 16'h200;
			16'h33e9: y = 16'h200;
			16'h33ea: y = 16'h200;
			16'h33eb: y = 16'h200;
			16'h33ec: y = 16'h200;
			16'h33ed: y = 16'h200;
			16'h33ee: y = 16'h200;
			16'h33ef: y = 16'h200;
			16'h33f0: y = 16'h200;
			16'h33f1: y = 16'h200;
			16'h33f2: y = 16'h200;
			16'h33f3: y = 16'h200;
			16'h33f4: y = 16'h200;
			16'h33f5: y = 16'h200;
			16'h33f6: y = 16'h200;
			16'h33f7: y = 16'h200;
			16'h33f8: y = 16'h200;
			16'h33f9: y = 16'h200;
			16'h33fa: y = 16'h200;
			16'h33fb: y = 16'h200;
			16'h33fc: y = 16'h200;
			16'h33fd: y = 16'h200;
			16'h33fe: y = 16'h200;
			16'h33ff: y = 16'h200;
			16'h3400: y = 16'h200;
			16'h3401: y = 16'h200;
			16'h3402: y = 16'h200;
			16'h3403: y = 16'h200;
			16'h3404: y = 16'h200;
			16'h3405: y = 16'h200;
			16'h3406: y = 16'h200;
			16'h3407: y = 16'h200;
			16'h3408: y = 16'h200;
			16'h3409: y = 16'h200;
			16'h340a: y = 16'h200;
			16'h340b: y = 16'h200;
			16'h340c: y = 16'h200;
			16'h340d: y = 16'h200;
			16'h340e: y = 16'h200;
			16'h340f: y = 16'h200;
			16'h3410: y = 16'h200;
			16'h3411: y = 16'h200;
			16'h3412: y = 16'h200;
			16'h3413: y = 16'h200;
			16'h3414: y = 16'h200;
			16'h3415: y = 16'h200;
			16'h3416: y = 16'h200;
			16'h3417: y = 16'h200;
			16'h3418: y = 16'h200;
			16'h3419: y = 16'h200;
			16'h341a: y = 16'h200;
			16'h341b: y = 16'h200;
			16'h341c: y = 16'h200;
			16'h341d: y = 16'h200;
			16'h341e: y = 16'h200;
			16'h341f: y = 16'h200;
			16'h3420: y = 16'h200;
			16'h3421: y = 16'h200;
			16'h3422: y = 16'h200;
			16'h3423: y = 16'h200;
			16'h3424: y = 16'h200;
			16'h3425: y = 16'h200;
			16'h3426: y = 16'h200;
			16'h3427: y = 16'h200;
			16'h3428: y = 16'h200;
			16'h3429: y = 16'h200;
			16'h342a: y = 16'h200;
			16'h342b: y = 16'h200;
			16'h342c: y = 16'h200;
			16'h342d: y = 16'h200;
			16'h342e: y = 16'h200;
			16'h342f: y = 16'h200;
			16'h3430: y = 16'h200;
			16'h3431: y = 16'h200;
			16'h3432: y = 16'h200;
			16'h3433: y = 16'h200;
			16'h3434: y = 16'h200;
			16'h3435: y = 16'h200;
			16'h3436: y = 16'h200;
			16'h3437: y = 16'h200;
			16'h3438: y = 16'h200;
			16'h3439: y = 16'h200;
			16'h343a: y = 16'h200;
			16'h343b: y = 16'h200;
			16'h343c: y = 16'h200;
			16'h343d: y = 16'h200;
			16'h343e: y = 16'h200;
			16'h343f: y = 16'h200;
			16'h3440: y = 16'h200;
			16'h3441: y = 16'h200;
			16'h3442: y = 16'h200;
			16'h3443: y = 16'h200;
			16'h3444: y = 16'h200;
			16'h3445: y = 16'h200;
			16'h3446: y = 16'h200;
			16'h3447: y = 16'h200;
			16'h3448: y = 16'h200;
			16'h3449: y = 16'h200;
			16'h344a: y = 16'h200;
			16'h344b: y = 16'h200;
			16'h344c: y = 16'h200;
			16'h344d: y = 16'h200;
			16'h344e: y = 16'h200;
			16'h344f: y = 16'h200;
			16'h3450: y = 16'h200;
			16'h3451: y = 16'h200;
			16'h3452: y = 16'h200;
			16'h3453: y = 16'h200;
			16'h3454: y = 16'h200;
			16'h3455: y = 16'h200;
			16'h3456: y = 16'h200;
			16'h3457: y = 16'h200;
			16'h3458: y = 16'h200;
			16'h3459: y = 16'h200;
			16'h345a: y = 16'h200;
			16'h345b: y = 16'h200;
			16'h345c: y = 16'h200;
			16'h345d: y = 16'h200;
			16'h345e: y = 16'h200;
			16'h345f: y = 16'h200;
			16'h3460: y = 16'h200;
			16'h3461: y = 16'h200;
			16'h3462: y = 16'h200;
			16'h3463: y = 16'h200;
			16'h3464: y = 16'h200;
			16'h3465: y = 16'h200;
			16'h3466: y = 16'h200;
			16'h3467: y = 16'h200;
			16'h3468: y = 16'h200;
			16'h3469: y = 16'h200;
			16'h346a: y = 16'h200;
			16'h346b: y = 16'h200;
			16'h346c: y = 16'h200;
			16'h346d: y = 16'h200;
			16'h346e: y = 16'h200;
			16'h346f: y = 16'h200;
			16'h3470: y = 16'h200;
			16'h3471: y = 16'h200;
			16'h3472: y = 16'h200;
			16'h3473: y = 16'h200;
			16'h3474: y = 16'h200;
			16'h3475: y = 16'h200;
			16'h3476: y = 16'h200;
			16'h3477: y = 16'h200;
			16'h3478: y = 16'h200;
			16'h3479: y = 16'h200;
			16'h347a: y = 16'h200;
			16'h347b: y = 16'h200;
			16'h347c: y = 16'h200;
			16'h347d: y = 16'h200;
			16'h347e: y = 16'h200;
			16'h347f: y = 16'h200;
			16'h3480: y = 16'h200;
			16'h3481: y = 16'h200;
			16'h3482: y = 16'h200;
			16'h3483: y = 16'h200;
			16'h3484: y = 16'h200;
			16'h3485: y = 16'h200;
			16'h3486: y = 16'h200;
			16'h3487: y = 16'h200;
			16'h3488: y = 16'h200;
			16'h3489: y = 16'h200;
			16'h348a: y = 16'h200;
			16'h348b: y = 16'h200;
			16'h348c: y = 16'h200;
			16'h348d: y = 16'h200;
			16'h348e: y = 16'h200;
			16'h348f: y = 16'h200;
			16'h3490: y = 16'h200;
			16'h3491: y = 16'h200;
			16'h3492: y = 16'h200;
			16'h3493: y = 16'h200;
			16'h3494: y = 16'h200;
			16'h3495: y = 16'h200;
			16'h3496: y = 16'h200;
			16'h3497: y = 16'h200;
			16'h3498: y = 16'h200;
			16'h3499: y = 16'h200;
			16'h349a: y = 16'h200;
			16'h349b: y = 16'h200;
			16'h349c: y = 16'h200;
			16'h349d: y = 16'h200;
			16'h349e: y = 16'h200;
			16'h349f: y = 16'h200;
			16'h34a0: y = 16'h200;
			16'h34a1: y = 16'h200;
			16'h34a2: y = 16'h200;
			16'h34a3: y = 16'h200;
			16'h34a4: y = 16'h200;
			16'h34a5: y = 16'h200;
			16'h34a6: y = 16'h200;
			16'h34a7: y = 16'h200;
			16'h34a8: y = 16'h200;
			16'h34a9: y = 16'h200;
			16'h34aa: y = 16'h200;
			16'h34ab: y = 16'h200;
			16'h34ac: y = 16'h200;
			16'h34ad: y = 16'h200;
			16'h34ae: y = 16'h200;
			16'h34af: y = 16'h200;
			16'h34b0: y = 16'h200;
			16'h34b1: y = 16'h200;
			16'h34b2: y = 16'h200;
			16'h34b3: y = 16'h200;
			16'h34b4: y = 16'h200;
			16'h34b5: y = 16'h200;
			16'h34b6: y = 16'h200;
			16'h34b7: y = 16'h200;
			16'h34b8: y = 16'h200;
			16'h34b9: y = 16'h200;
			16'h34ba: y = 16'h200;
			16'h34bb: y = 16'h200;
			16'h34bc: y = 16'h200;
			16'h34bd: y = 16'h200;
			16'h34be: y = 16'h200;
			16'h34bf: y = 16'h200;
			16'h34c0: y = 16'h200;
			16'h34c1: y = 16'h200;
			16'h34c2: y = 16'h200;
			16'h34c3: y = 16'h200;
			16'h34c4: y = 16'h200;
			16'h34c5: y = 16'h200;
			16'h34c6: y = 16'h200;
			16'h34c7: y = 16'h200;
			16'h34c8: y = 16'h200;
			16'h34c9: y = 16'h200;
			16'h34ca: y = 16'h200;
			16'h34cb: y = 16'h200;
			16'h34cc: y = 16'h200;
			16'h34cd: y = 16'h200;
			16'h34ce: y = 16'h200;
			16'h34cf: y = 16'h200;
			16'h34d0: y = 16'h200;
			16'h34d1: y = 16'h200;
			16'h34d2: y = 16'h200;
			16'h34d3: y = 16'h200;
			16'h34d4: y = 16'h200;
			16'h34d5: y = 16'h200;
			16'h34d6: y = 16'h200;
			16'h34d7: y = 16'h200;
			16'h34d8: y = 16'h200;
			16'h34d9: y = 16'h200;
			16'h34da: y = 16'h200;
			16'h34db: y = 16'h200;
			16'h34dc: y = 16'h200;
			16'h34dd: y = 16'h200;
			16'h34de: y = 16'h200;
			16'h34df: y = 16'h200;
			16'h34e0: y = 16'h200;
			16'h34e1: y = 16'h200;
			16'h34e2: y = 16'h200;
			16'h34e3: y = 16'h200;
			16'h34e4: y = 16'h200;
			16'h34e5: y = 16'h200;
			16'h34e6: y = 16'h200;
			16'h34e7: y = 16'h200;
			16'h34e8: y = 16'h200;
			16'h34e9: y = 16'h200;
			16'h34ea: y = 16'h200;
			16'h34eb: y = 16'h200;
			16'h34ec: y = 16'h200;
			16'h34ed: y = 16'h200;
			16'h34ee: y = 16'h200;
			16'h34ef: y = 16'h200;
			16'h34f0: y = 16'h200;
			16'h34f1: y = 16'h200;
			16'h34f2: y = 16'h200;
			16'h34f3: y = 16'h200;
			16'h34f4: y = 16'h200;
			16'h34f5: y = 16'h200;
			16'h34f6: y = 16'h200;
			16'h34f7: y = 16'h200;
			16'h34f8: y = 16'h200;
			16'h34f9: y = 16'h200;
			16'h34fa: y = 16'h200;
			16'h34fb: y = 16'h200;
			16'h34fc: y = 16'h200;
			16'h34fd: y = 16'h200;
			16'h34fe: y = 16'h200;
			16'h34ff: y = 16'h200;
			16'h3500: y = 16'h200;
			16'h3501: y = 16'h200;
			16'h3502: y = 16'h200;
			16'h3503: y = 16'h200;
			16'h3504: y = 16'h200;
			16'h3505: y = 16'h200;
			16'h3506: y = 16'h200;
			16'h3507: y = 16'h200;
			16'h3508: y = 16'h200;
			16'h3509: y = 16'h200;
			16'h350a: y = 16'h200;
			16'h350b: y = 16'h200;
			16'h350c: y = 16'h200;
			16'h350d: y = 16'h200;
			16'h350e: y = 16'h200;
			16'h350f: y = 16'h200;
			16'h3510: y = 16'h200;
			16'h3511: y = 16'h200;
			16'h3512: y = 16'h200;
			16'h3513: y = 16'h200;
			16'h3514: y = 16'h200;
			16'h3515: y = 16'h200;
			16'h3516: y = 16'h200;
			16'h3517: y = 16'h200;
			16'h3518: y = 16'h200;
			16'h3519: y = 16'h200;
			16'h351a: y = 16'h200;
			16'h351b: y = 16'h200;
			16'h351c: y = 16'h200;
			16'h351d: y = 16'h200;
			16'h351e: y = 16'h200;
			16'h351f: y = 16'h200;
			16'h3520: y = 16'h200;
			16'h3521: y = 16'h200;
			16'h3522: y = 16'h200;
			16'h3523: y = 16'h200;
			16'h3524: y = 16'h200;
			16'h3525: y = 16'h200;
			16'h3526: y = 16'h200;
			16'h3527: y = 16'h200;
			16'h3528: y = 16'h200;
			16'h3529: y = 16'h200;
			16'h352a: y = 16'h200;
			16'h352b: y = 16'h200;
			16'h352c: y = 16'h200;
			16'h352d: y = 16'h200;
			16'h352e: y = 16'h200;
			16'h352f: y = 16'h200;
			16'h3530: y = 16'h200;
			16'h3531: y = 16'h200;
			16'h3532: y = 16'h200;
			16'h3533: y = 16'h200;
			16'h3534: y = 16'h200;
			16'h3535: y = 16'h200;
			16'h3536: y = 16'h200;
			16'h3537: y = 16'h200;
			16'h3538: y = 16'h200;
			16'h3539: y = 16'h200;
			16'h353a: y = 16'h200;
			16'h353b: y = 16'h200;
			16'h353c: y = 16'h200;
			16'h353d: y = 16'h200;
			16'h353e: y = 16'h200;
			16'h353f: y = 16'h200;
			16'h3540: y = 16'h200;
			16'h3541: y = 16'h200;
			16'h3542: y = 16'h200;
			16'h3543: y = 16'h200;
			16'h3544: y = 16'h200;
			16'h3545: y = 16'h200;
			16'h3546: y = 16'h200;
			16'h3547: y = 16'h200;
			16'h3548: y = 16'h200;
			16'h3549: y = 16'h200;
			16'h354a: y = 16'h200;
			16'h354b: y = 16'h200;
			16'h354c: y = 16'h200;
			16'h354d: y = 16'h200;
			16'h354e: y = 16'h200;
			16'h354f: y = 16'h200;
			16'h3550: y = 16'h200;
			16'h3551: y = 16'h200;
			16'h3552: y = 16'h200;
			16'h3553: y = 16'h200;
			16'h3554: y = 16'h200;
			16'h3555: y = 16'h200;
			16'h3556: y = 16'h200;
			16'h3557: y = 16'h200;
			16'h3558: y = 16'h200;
			16'h3559: y = 16'h200;
			16'h355a: y = 16'h200;
			16'h355b: y = 16'h200;
			16'h355c: y = 16'h200;
			16'h355d: y = 16'h200;
			16'h355e: y = 16'h200;
			16'h355f: y = 16'h200;
			16'h3560: y = 16'h200;
			16'h3561: y = 16'h200;
			16'h3562: y = 16'h200;
			16'h3563: y = 16'h200;
			16'h3564: y = 16'h200;
			16'h3565: y = 16'h200;
			16'h3566: y = 16'h200;
			16'h3567: y = 16'h200;
			16'h3568: y = 16'h200;
			16'h3569: y = 16'h200;
			16'h356a: y = 16'h200;
			16'h356b: y = 16'h200;
			16'h356c: y = 16'h200;
			16'h356d: y = 16'h200;
			16'h356e: y = 16'h200;
			16'h356f: y = 16'h200;
			16'h3570: y = 16'h200;
			16'h3571: y = 16'h200;
			16'h3572: y = 16'h200;
			16'h3573: y = 16'h200;
			16'h3574: y = 16'h200;
			16'h3575: y = 16'h200;
			16'h3576: y = 16'h200;
			16'h3577: y = 16'h200;
			16'h3578: y = 16'h200;
			16'h3579: y = 16'h200;
			16'h357a: y = 16'h200;
			16'h357b: y = 16'h200;
			16'h357c: y = 16'h200;
			16'h357d: y = 16'h200;
			16'h357e: y = 16'h200;
			16'h357f: y = 16'h200;
			16'h3580: y = 16'h200;
			16'h3581: y = 16'h200;
			16'h3582: y = 16'h200;
			16'h3583: y = 16'h200;
			16'h3584: y = 16'h200;
			16'h3585: y = 16'h200;
			16'h3586: y = 16'h200;
			16'h3587: y = 16'h200;
			16'h3588: y = 16'h200;
			16'h3589: y = 16'h200;
			16'h358a: y = 16'h200;
			16'h358b: y = 16'h200;
			16'h358c: y = 16'h200;
			16'h358d: y = 16'h200;
			16'h358e: y = 16'h200;
			16'h358f: y = 16'h200;
			16'h3590: y = 16'h200;
			16'h3591: y = 16'h200;
			16'h3592: y = 16'h200;
			16'h3593: y = 16'h200;
			16'h3594: y = 16'h200;
			16'h3595: y = 16'h200;
			16'h3596: y = 16'h200;
			16'h3597: y = 16'h200;
			16'h3598: y = 16'h200;
			16'h3599: y = 16'h200;
			16'h359a: y = 16'h200;
			16'h359b: y = 16'h200;
			16'h359c: y = 16'h200;
			16'h359d: y = 16'h200;
			16'h359e: y = 16'h200;
			16'h359f: y = 16'h200;
			16'h35a0: y = 16'h200;
			16'h35a1: y = 16'h200;
			16'h35a2: y = 16'h200;
			16'h35a3: y = 16'h200;
			16'h35a4: y = 16'h200;
			16'h35a5: y = 16'h200;
			16'h35a6: y = 16'h200;
			16'h35a7: y = 16'h200;
			16'h35a8: y = 16'h200;
			16'h35a9: y = 16'h200;
			16'h35aa: y = 16'h200;
			16'h35ab: y = 16'h200;
			16'h35ac: y = 16'h200;
			16'h35ad: y = 16'h200;
			16'h35ae: y = 16'h200;
			16'h35af: y = 16'h200;
			16'h35b0: y = 16'h200;
			16'h35b1: y = 16'h200;
			16'h35b2: y = 16'h200;
			16'h35b3: y = 16'h200;
			16'h35b4: y = 16'h200;
			16'h35b5: y = 16'h200;
			16'h35b6: y = 16'h200;
			16'h35b7: y = 16'h200;
			16'h35b8: y = 16'h200;
			16'h35b9: y = 16'h200;
			16'h35ba: y = 16'h200;
			16'h35bb: y = 16'h200;
			16'h35bc: y = 16'h200;
			16'h35bd: y = 16'h200;
			16'h35be: y = 16'h200;
			16'h35bf: y = 16'h200;
			16'h35c0: y = 16'h200;
			16'h35c1: y = 16'h200;
			16'h35c2: y = 16'h200;
			16'h35c3: y = 16'h200;
			16'h35c4: y = 16'h200;
			16'h35c5: y = 16'h200;
			16'h35c6: y = 16'h200;
			16'h35c7: y = 16'h200;
			16'h35c8: y = 16'h200;
			16'h35c9: y = 16'h200;
			16'h35ca: y = 16'h200;
			16'h35cb: y = 16'h200;
			16'h35cc: y = 16'h200;
			16'h35cd: y = 16'h200;
			16'h35ce: y = 16'h200;
			16'h35cf: y = 16'h200;
			16'h35d0: y = 16'h200;
			16'h35d1: y = 16'h200;
			16'h35d2: y = 16'h200;
			16'h35d3: y = 16'h200;
			16'h35d4: y = 16'h200;
			16'h35d5: y = 16'h200;
			16'h35d6: y = 16'h200;
			16'h35d7: y = 16'h200;
			16'h35d8: y = 16'h200;
			16'h35d9: y = 16'h200;
			16'h35da: y = 16'h200;
			16'h35db: y = 16'h200;
			16'h35dc: y = 16'h200;
			16'h35dd: y = 16'h200;
			16'h35de: y = 16'h200;
			16'h35df: y = 16'h200;
			16'h35e0: y = 16'h200;
			16'h35e1: y = 16'h200;
			16'h35e2: y = 16'h200;
			16'h35e3: y = 16'h200;
			16'h35e4: y = 16'h200;
			16'h35e5: y = 16'h200;
			16'h35e6: y = 16'h200;
			16'h35e7: y = 16'h200;
			16'h35e8: y = 16'h200;
			16'h35e9: y = 16'h200;
			16'h35ea: y = 16'h200;
			16'h35eb: y = 16'h200;
			16'h35ec: y = 16'h200;
			16'h35ed: y = 16'h200;
			16'h35ee: y = 16'h200;
			16'h35ef: y = 16'h200;
			16'h35f0: y = 16'h200;
			16'h35f1: y = 16'h200;
			16'h35f2: y = 16'h200;
			16'h35f3: y = 16'h200;
			16'h35f4: y = 16'h200;
			16'h35f5: y = 16'h200;
			16'h35f6: y = 16'h200;
			16'h35f7: y = 16'h200;
			16'h35f8: y = 16'h200;
			16'h35f9: y = 16'h200;
			16'h35fa: y = 16'h200;
			16'h35fb: y = 16'h200;
			16'h35fc: y = 16'h200;
			16'h35fd: y = 16'h200;
			16'h35fe: y = 16'h200;
			16'h35ff: y = 16'h200;
			16'h3600: y = 16'h200;
			16'h3601: y = 16'h200;
			16'h3602: y = 16'h200;
			16'h3603: y = 16'h200;
			16'h3604: y = 16'h200;
			16'h3605: y = 16'h200;
			16'h3606: y = 16'h200;
			16'h3607: y = 16'h200;
			16'h3608: y = 16'h200;
			16'h3609: y = 16'h200;
			16'h360a: y = 16'h200;
			16'h360b: y = 16'h200;
			16'h360c: y = 16'h200;
			16'h360d: y = 16'h200;
			16'h360e: y = 16'h200;
			16'h360f: y = 16'h200;
			16'h3610: y = 16'h200;
			16'h3611: y = 16'h200;
			16'h3612: y = 16'h200;
			16'h3613: y = 16'h200;
			16'h3614: y = 16'h200;
			16'h3615: y = 16'h200;
			16'h3616: y = 16'h200;
			16'h3617: y = 16'h200;
			16'h3618: y = 16'h200;
			16'h3619: y = 16'h200;
			16'h361a: y = 16'h200;
			16'h361b: y = 16'h200;
			16'h361c: y = 16'h200;
			16'h361d: y = 16'h200;
			16'h361e: y = 16'h200;
			16'h361f: y = 16'h200;
			16'h3620: y = 16'h200;
			16'h3621: y = 16'h200;
			16'h3622: y = 16'h200;
			16'h3623: y = 16'h200;
			16'h3624: y = 16'h200;
			16'h3625: y = 16'h200;
			16'h3626: y = 16'h200;
			16'h3627: y = 16'h200;
			16'h3628: y = 16'h200;
			16'h3629: y = 16'h200;
			16'h362a: y = 16'h200;
			16'h362b: y = 16'h200;
			16'h362c: y = 16'h200;
			16'h362d: y = 16'h200;
			16'h362e: y = 16'h200;
			16'h362f: y = 16'h200;
			16'h3630: y = 16'h200;
			16'h3631: y = 16'h200;
			16'h3632: y = 16'h200;
			16'h3633: y = 16'h200;
			16'h3634: y = 16'h200;
			16'h3635: y = 16'h200;
			16'h3636: y = 16'h200;
			16'h3637: y = 16'h200;
			16'h3638: y = 16'h200;
			16'h3639: y = 16'h200;
			16'h363a: y = 16'h200;
			16'h363b: y = 16'h200;
			16'h363c: y = 16'h200;
			16'h363d: y = 16'h200;
			16'h363e: y = 16'h200;
			16'h363f: y = 16'h200;
			16'h3640: y = 16'h200;
			16'h3641: y = 16'h200;
			16'h3642: y = 16'h200;
			16'h3643: y = 16'h200;
			16'h3644: y = 16'h200;
			16'h3645: y = 16'h200;
			16'h3646: y = 16'h200;
			16'h3647: y = 16'h200;
			16'h3648: y = 16'h200;
			16'h3649: y = 16'h200;
			16'h364a: y = 16'h200;
			16'h364b: y = 16'h200;
			16'h364c: y = 16'h200;
			16'h364d: y = 16'h200;
			16'h364e: y = 16'h200;
			16'h364f: y = 16'h200;
			16'h3650: y = 16'h200;
			16'h3651: y = 16'h200;
			16'h3652: y = 16'h200;
			16'h3653: y = 16'h200;
			16'h3654: y = 16'h200;
			16'h3655: y = 16'h200;
			16'h3656: y = 16'h200;
			16'h3657: y = 16'h200;
			16'h3658: y = 16'h200;
			16'h3659: y = 16'h200;
			16'h365a: y = 16'h200;
			16'h365b: y = 16'h200;
			16'h365c: y = 16'h200;
			16'h365d: y = 16'h200;
			16'h365e: y = 16'h200;
			16'h365f: y = 16'h200;
			16'h3660: y = 16'h200;
			16'h3661: y = 16'h200;
			16'h3662: y = 16'h200;
			16'h3663: y = 16'h200;
			16'h3664: y = 16'h200;
			16'h3665: y = 16'h200;
			16'h3666: y = 16'h200;
			16'h3667: y = 16'h200;
			16'h3668: y = 16'h200;
			16'h3669: y = 16'h200;
			16'h366a: y = 16'h200;
			16'h366b: y = 16'h200;
			16'h366c: y = 16'h200;
			16'h366d: y = 16'h200;
			16'h366e: y = 16'h200;
			16'h366f: y = 16'h200;
			16'h3670: y = 16'h200;
			16'h3671: y = 16'h200;
			16'h3672: y = 16'h200;
			16'h3673: y = 16'h200;
			16'h3674: y = 16'h200;
			16'h3675: y = 16'h200;
			16'h3676: y = 16'h200;
			16'h3677: y = 16'h200;
			16'h3678: y = 16'h200;
			16'h3679: y = 16'h200;
			16'h367a: y = 16'h200;
			16'h367b: y = 16'h200;
			16'h367c: y = 16'h200;
			16'h367d: y = 16'h200;
			16'h367e: y = 16'h200;
			16'h367f: y = 16'h200;
			16'h3680: y = 16'h200;
			16'h3681: y = 16'h200;
			16'h3682: y = 16'h200;
			16'h3683: y = 16'h200;
			16'h3684: y = 16'h200;
			16'h3685: y = 16'h200;
			16'h3686: y = 16'h200;
			16'h3687: y = 16'h200;
			16'h3688: y = 16'h200;
			16'h3689: y = 16'h200;
			16'h368a: y = 16'h200;
			16'h368b: y = 16'h200;
			16'h368c: y = 16'h200;
			16'h368d: y = 16'h200;
			16'h368e: y = 16'h200;
			16'h368f: y = 16'h200;
			16'h3690: y = 16'h200;
			16'h3691: y = 16'h200;
			16'h3692: y = 16'h200;
			16'h3693: y = 16'h200;
			16'h3694: y = 16'h200;
			16'h3695: y = 16'h200;
			16'h3696: y = 16'h200;
			16'h3697: y = 16'h200;
			16'h3698: y = 16'h200;
			16'h3699: y = 16'h200;
			16'h369a: y = 16'h200;
			16'h369b: y = 16'h200;
			16'h369c: y = 16'h200;
			16'h369d: y = 16'h200;
			16'h369e: y = 16'h200;
			16'h369f: y = 16'h200;
			16'h36a0: y = 16'h200;
			16'h36a1: y = 16'h200;
			16'h36a2: y = 16'h200;
			16'h36a3: y = 16'h200;
			16'h36a4: y = 16'h200;
			16'h36a5: y = 16'h200;
			16'h36a6: y = 16'h200;
			16'h36a7: y = 16'h200;
			16'h36a8: y = 16'h200;
			16'h36a9: y = 16'h200;
			16'h36aa: y = 16'h200;
			16'h36ab: y = 16'h200;
			16'h36ac: y = 16'h200;
			16'h36ad: y = 16'h200;
			16'h36ae: y = 16'h200;
			16'h36af: y = 16'h200;
			16'h36b0: y = 16'h200;
			16'h36b1: y = 16'h200;
			16'h36b2: y = 16'h200;
			16'h36b3: y = 16'h200;
			16'h36b4: y = 16'h200;
			16'h36b5: y = 16'h200;
			16'h36b6: y = 16'h200;
			16'h36b7: y = 16'h200;
			16'h36b8: y = 16'h200;
			16'h36b9: y = 16'h200;
			16'h36ba: y = 16'h200;
			16'h36bb: y = 16'h200;
			16'h36bc: y = 16'h200;
			16'h36bd: y = 16'h200;
			16'h36be: y = 16'h200;
			16'h36bf: y = 16'h200;
			16'h36c0: y = 16'h200;
			16'h36c1: y = 16'h200;
			16'h36c2: y = 16'h200;
			16'h36c3: y = 16'h200;
			16'h36c4: y = 16'h200;
			16'h36c5: y = 16'h200;
			16'h36c6: y = 16'h200;
			16'h36c7: y = 16'h200;
			16'h36c8: y = 16'h200;
			16'h36c9: y = 16'h200;
			16'h36ca: y = 16'h200;
			16'h36cb: y = 16'h200;
			16'h36cc: y = 16'h200;
			16'h36cd: y = 16'h200;
			16'h36ce: y = 16'h200;
			16'h36cf: y = 16'h200;
			16'h36d0: y = 16'h200;
			16'h36d1: y = 16'h200;
			16'h36d2: y = 16'h200;
			16'h36d3: y = 16'h200;
			16'h36d4: y = 16'h200;
			16'h36d5: y = 16'h200;
			16'h36d6: y = 16'h200;
			16'h36d7: y = 16'h200;
			16'h36d8: y = 16'h200;
			16'h36d9: y = 16'h200;
			16'h36da: y = 16'h200;
			16'h36db: y = 16'h200;
			16'h36dc: y = 16'h200;
			16'h36dd: y = 16'h200;
			16'h36de: y = 16'h200;
			16'h36df: y = 16'h200;
			16'h36e0: y = 16'h200;
			16'h36e1: y = 16'h200;
			16'h36e2: y = 16'h200;
			16'h36e3: y = 16'h200;
			16'h36e4: y = 16'h200;
			16'h36e5: y = 16'h200;
			16'h36e6: y = 16'h200;
			16'h36e7: y = 16'h200;
			16'h36e8: y = 16'h200;
			16'h36e9: y = 16'h200;
			16'h36ea: y = 16'h200;
			16'h36eb: y = 16'h200;
			16'h36ec: y = 16'h200;
			16'h36ed: y = 16'h200;
			16'h36ee: y = 16'h200;
			16'h36ef: y = 16'h200;
			16'h36f0: y = 16'h200;
			16'h36f1: y = 16'h200;
			16'h36f2: y = 16'h200;
			16'h36f3: y = 16'h200;
			16'h36f4: y = 16'h200;
			16'h36f5: y = 16'h200;
			16'h36f6: y = 16'h200;
			16'h36f7: y = 16'h200;
			16'h36f8: y = 16'h200;
			16'h36f9: y = 16'h200;
			16'h36fa: y = 16'h200;
			16'h36fb: y = 16'h200;
			16'h36fc: y = 16'h200;
			16'h36fd: y = 16'h200;
			16'h36fe: y = 16'h200;
			16'h36ff: y = 16'h200;
			16'h3700: y = 16'h200;
			16'h3701: y = 16'h200;
			16'h3702: y = 16'h200;
			16'h3703: y = 16'h200;
			16'h3704: y = 16'h200;
			16'h3705: y = 16'h200;
			16'h3706: y = 16'h200;
			16'h3707: y = 16'h200;
			16'h3708: y = 16'h200;
			16'h3709: y = 16'h200;
			16'h370a: y = 16'h200;
			16'h370b: y = 16'h200;
			16'h370c: y = 16'h200;
			16'h370d: y = 16'h200;
			16'h370e: y = 16'h200;
			16'h370f: y = 16'h200;
			16'h3710: y = 16'h200;
			16'h3711: y = 16'h200;
			16'h3712: y = 16'h200;
			16'h3713: y = 16'h200;
			16'h3714: y = 16'h200;
			16'h3715: y = 16'h200;
			16'h3716: y = 16'h200;
			16'h3717: y = 16'h200;
			16'h3718: y = 16'h200;
			16'h3719: y = 16'h200;
			16'h371a: y = 16'h200;
			16'h371b: y = 16'h200;
			16'h371c: y = 16'h200;
			16'h371d: y = 16'h200;
			16'h371e: y = 16'h200;
			16'h371f: y = 16'h200;
			16'h3720: y = 16'h200;
			16'h3721: y = 16'h200;
			16'h3722: y = 16'h200;
			16'h3723: y = 16'h200;
			16'h3724: y = 16'h200;
			16'h3725: y = 16'h200;
			16'h3726: y = 16'h200;
			16'h3727: y = 16'h200;
			16'h3728: y = 16'h200;
			16'h3729: y = 16'h200;
			16'h372a: y = 16'h200;
			16'h372b: y = 16'h200;
			16'h372c: y = 16'h200;
			16'h372d: y = 16'h200;
			16'h372e: y = 16'h200;
			16'h372f: y = 16'h200;
			16'h3730: y = 16'h200;
			16'h3731: y = 16'h200;
			16'h3732: y = 16'h200;
			16'h3733: y = 16'h200;
			16'h3734: y = 16'h200;
			16'h3735: y = 16'h200;
			16'h3736: y = 16'h200;
			16'h3737: y = 16'h200;
			16'h3738: y = 16'h200;
			16'h3739: y = 16'h200;
			16'h373a: y = 16'h200;
			16'h373b: y = 16'h200;
			16'h373c: y = 16'h200;
			16'h373d: y = 16'h200;
			16'h373e: y = 16'h200;
			16'h373f: y = 16'h200;
			16'h3740: y = 16'h200;
			16'h3741: y = 16'h200;
			16'h3742: y = 16'h200;
			16'h3743: y = 16'h200;
			16'h3744: y = 16'h200;
			16'h3745: y = 16'h200;
			16'h3746: y = 16'h200;
			16'h3747: y = 16'h200;
			16'h3748: y = 16'h200;
			16'h3749: y = 16'h200;
			16'h374a: y = 16'h200;
			16'h374b: y = 16'h200;
			16'h374c: y = 16'h200;
			16'h374d: y = 16'h200;
			16'h374e: y = 16'h200;
			16'h374f: y = 16'h200;
			16'h3750: y = 16'h200;
			16'h3751: y = 16'h200;
			16'h3752: y = 16'h200;
			16'h3753: y = 16'h200;
			16'h3754: y = 16'h200;
			16'h3755: y = 16'h200;
			16'h3756: y = 16'h200;
			16'h3757: y = 16'h200;
			16'h3758: y = 16'h200;
			16'h3759: y = 16'h200;
			16'h375a: y = 16'h200;
			16'h375b: y = 16'h200;
			16'h375c: y = 16'h200;
			16'h375d: y = 16'h200;
			16'h375e: y = 16'h200;
			16'h375f: y = 16'h200;
			16'h3760: y = 16'h200;
			16'h3761: y = 16'h200;
			16'h3762: y = 16'h200;
			16'h3763: y = 16'h200;
			16'h3764: y = 16'h200;
			16'h3765: y = 16'h200;
			16'h3766: y = 16'h200;
			16'h3767: y = 16'h200;
			16'h3768: y = 16'h200;
			16'h3769: y = 16'h200;
			16'h376a: y = 16'h200;
			16'h376b: y = 16'h200;
			16'h376c: y = 16'h200;
			16'h376d: y = 16'h200;
			16'h376e: y = 16'h200;
			16'h376f: y = 16'h200;
			16'h3770: y = 16'h200;
			16'h3771: y = 16'h200;
			16'h3772: y = 16'h200;
			16'h3773: y = 16'h200;
			16'h3774: y = 16'h200;
			16'h3775: y = 16'h200;
			16'h3776: y = 16'h200;
			16'h3777: y = 16'h200;
			16'h3778: y = 16'h200;
			16'h3779: y = 16'h200;
			16'h377a: y = 16'h200;
			16'h377b: y = 16'h200;
			16'h377c: y = 16'h200;
			16'h377d: y = 16'h200;
			16'h377e: y = 16'h200;
			16'h377f: y = 16'h200;
			16'h3780: y = 16'h200;
			16'h3781: y = 16'h200;
			16'h3782: y = 16'h200;
			16'h3783: y = 16'h200;
			16'h3784: y = 16'h200;
			16'h3785: y = 16'h200;
			16'h3786: y = 16'h200;
			16'h3787: y = 16'h200;
			16'h3788: y = 16'h200;
			16'h3789: y = 16'h200;
			16'h378a: y = 16'h200;
			16'h378b: y = 16'h200;
			16'h378c: y = 16'h200;
			16'h378d: y = 16'h200;
			16'h378e: y = 16'h200;
			16'h378f: y = 16'h200;
			16'h3790: y = 16'h200;
			16'h3791: y = 16'h200;
			16'h3792: y = 16'h200;
			16'h3793: y = 16'h200;
			16'h3794: y = 16'h200;
			16'h3795: y = 16'h200;
			16'h3796: y = 16'h200;
			16'h3797: y = 16'h200;
			16'h3798: y = 16'h200;
			16'h3799: y = 16'h200;
			16'h379a: y = 16'h200;
			16'h379b: y = 16'h200;
			16'h379c: y = 16'h200;
			16'h379d: y = 16'h200;
			16'h379e: y = 16'h200;
			16'h379f: y = 16'h200;
			16'h37a0: y = 16'h200;
			16'h37a1: y = 16'h200;
			16'h37a2: y = 16'h200;
			16'h37a3: y = 16'h200;
			16'h37a4: y = 16'h200;
			16'h37a5: y = 16'h200;
			16'h37a6: y = 16'h200;
			16'h37a7: y = 16'h200;
			16'h37a8: y = 16'h200;
			16'h37a9: y = 16'h200;
			16'h37aa: y = 16'h200;
			16'h37ab: y = 16'h200;
			16'h37ac: y = 16'h200;
			16'h37ad: y = 16'h200;
			16'h37ae: y = 16'h200;
			16'h37af: y = 16'h200;
			16'h37b0: y = 16'h200;
			16'h37b1: y = 16'h200;
			16'h37b2: y = 16'h200;
			16'h37b3: y = 16'h200;
			16'h37b4: y = 16'h200;
			16'h37b5: y = 16'h200;
			16'h37b6: y = 16'h200;
			16'h37b7: y = 16'h200;
			16'h37b8: y = 16'h200;
			16'h37b9: y = 16'h200;
			16'h37ba: y = 16'h200;
			16'h37bb: y = 16'h200;
			16'h37bc: y = 16'h200;
			16'h37bd: y = 16'h200;
			16'h37be: y = 16'h200;
			16'h37bf: y = 16'h200;
			16'h37c0: y = 16'h200;
			16'h37c1: y = 16'h200;
			16'h37c2: y = 16'h200;
			16'h37c3: y = 16'h200;
			16'h37c4: y = 16'h200;
			16'h37c5: y = 16'h200;
			16'h37c6: y = 16'h200;
			16'h37c7: y = 16'h200;
			16'h37c8: y = 16'h200;
			16'h37c9: y = 16'h200;
			16'h37ca: y = 16'h200;
			16'h37cb: y = 16'h200;
			16'h37cc: y = 16'h200;
			16'h37cd: y = 16'h200;
			16'h37ce: y = 16'h200;
			16'h37cf: y = 16'h200;
			16'h37d0: y = 16'h200;
			16'h37d1: y = 16'h200;
			16'h37d2: y = 16'h200;
			16'h37d3: y = 16'h200;
			16'h37d4: y = 16'h200;
			16'h37d5: y = 16'h200;
			16'h37d6: y = 16'h200;
			16'h37d7: y = 16'h200;
			16'h37d8: y = 16'h200;
			16'h37d9: y = 16'h200;
			16'h37da: y = 16'h200;
			16'h37db: y = 16'h200;
			16'h37dc: y = 16'h200;
			16'h37dd: y = 16'h200;
			16'h37de: y = 16'h200;
			16'h37df: y = 16'h200;
			16'h37e0: y = 16'h200;
			16'h37e1: y = 16'h200;
			16'h37e2: y = 16'h200;
			16'h37e3: y = 16'h200;
			16'h37e4: y = 16'h200;
			16'h37e5: y = 16'h200;
			16'h37e6: y = 16'h200;
			16'h37e7: y = 16'h200;
			16'h37e8: y = 16'h200;
			16'h37e9: y = 16'h200;
			16'h37ea: y = 16'h200;
			16'h37eb: y = 16'h200;
			16'h37ec: y = 16'h200;
			16'h37ed: y = 16'h200;
			16'h37ee: y = 16'h200;
			16'h37ef: y = 16'h200;
			16'h37f0: y = 16'h200;
			16'h37f1: y = 16'h200;
			16'h37f2: y = 16'h200;
			16'h37f3: y = 16'h200;
			16'h37f4: y = 16'h200;
			16'h37f5: y = 16'h200;
			16'h37f6: y = 16'h200;
			16'h37f7: y = 16'h200;
			16'h37f8: y = 16'h200;
			16'h37f9: y = 16'h200;
			16'h37fa: y = 16'h200;
			16'h37fb: y = 16'h200;
			16'h37fc: y = 16'h200;
			16'h37fd: y = 16'h200;
			16'h37fe: y = 16'h200;
			16'h37ff: y = 16'h200;
			16'h3800: y = 16'h200;
			16'h3801: y = 16'h200;
			16'h3802: y = 16'h200;
			16'h3803: y = 16'h200;
			16'h3804: y = 16'h200;
			16'h3805: y = 16'h200;
			16'h3806: y = 16'h200;
			16'h3807: y = 16'h200;
			16'h3808: y = 16'h200;
			16'h3809: y = 16'h200;
			16'h380a: y = 16'h200;
			16'h380b: y = 16'h200;
			16'h380c: y = 16'h200;
			16'h380d: y = 16'h200;
			16'h380e: y = 16'h200;
			16'h380f: y = 16'h200;
			16'h3810: y = 16'h200;
			16'h3811: y = 16'h200;
			16'h3812: y = 16'h200;
			16'h3813: y = 16'h200;
			16'h3814: y = 16'h200;
			16'h3815: y = 16'h200;
			16'h3816: y = 16'h200;
			16'h3817: y = 16'h200;
			16'h3818: y = 16'h200;
			16'h3819: y = 16'h200;
			16'h381a: y = 16'h200;
			16'h381b: y = 16'h200;
			16'h381c: y = 16'h200;
			16'h381d: y = 16'h200;
			16'h381e: y = 16'h200;
			16'h381f: y = 16'h200;
			16'h3820: y = 16'h200;
			16'h3821: y = 16'h200;
			16'h3822: y = 16'h200;
			16'h3823: y = 16'h200;
			16'h3824: y = 16'h200;
			16'h3825: y = 16'h200;
			16'h3826: y = 16'h200;
			16'h3827: y = 16'h200;
			16'h3828: y = 16'h200;
			16'h3829: y = 16'h200;
			16'h382a: y = 16'h200;
			16'h382b: y = 16'h200;
			16'h382c: y = 16'h200;
			16'h382d: y = 16'h200;
			16'h382e: y = 16'h200;
			16'h382f: y = 16'h200;
			16'h3830: y = 16'h200;
			16'h3831: y = 16'h200;
			16'h3832: y = 16'h200;
			16'h3833: y = 16'h200;
			16'h3834: y = 16'h200;
			16'h3835: y = 16'h200;
			16'h3836: y = 16'h200;
			16'h3837: y = 16'h200;
			16'h3838: y = 16'h200;
			16'h3839: y = 16'h200;
			16'h383a: y = 16'h200;
			16'h383b: y = 16'h200;
			16'h383c: y = 16'h200;
			16'h383d: y = 16'h200;
			16'h383e: y = 16'h200;
			16'h383f: y = 16'h200;
			16'h3840: y = 16'h200;
			16'h3841: y = 16'h200;
			16'h3842: y = 16'h200;
			16'h3843: y = 16'h200;
			16'h3844: y = 16'h200;
			16'h3845: y = 16'h200;
			16'h3846: y = 16'h200;
			16'h3847: y = 16'h200;
			16'h3848: y = 16'h200;
			16'h3849: y = 16'h200;
			16'h384a: y = 16'h200;
			16'h384b: y = 16'h200;
			16'h384c: y = 16'h200;
			16'h384d: y = 16'h200;
			16'h384e: y = 16'h200;
			16'h384f: y = 16'h200;
			16'h3850: y = 16'h200;
			16'h3851: y = 16'h200;
			16'h3852: y = 16'h200;
			16'h3853: y = 16'h200;
			16'h3854: y = 16'h200;
			16'h3855: y = 16'h200;
			16'h3856: y = 16'h200;
			16'h3857: y = 16'h200;
			16'h3858: y = 16'h200;
			16'h3859: y = 16'h200;
			16'h385a: y = 16'h200;
			16'h385b: y = 16'h200;
			16'h385c: y = 16'h200;
			16'h385d: y = 16'h200;
			16'h385e: y = 16'h200;
			16'h385f: y = 16'h200;
			16'h3860: y = 16'h200;
			16'h3861: y = 16'h200;
			16'h3862: y = 16'h200;
			16'h3863: y = 16'h200;
			16'h3864: y = 16'h200;
			16'h3865: y = 16'h200;
			16'h3866: y = 16'h200;
			16'h3867: y = 16'h200;
			16'h3868: y = 16'h200;
			16'h3869: y = 16'h200;
			16'h386a: y = 16'h200;
			16'h386b: y = 16'h200;
			16'h386c: y = 16'h200;
			16'h386d: y = 16'h200;
			16'h386e: y = 16'h200;
			16'h386f: y = 16'h200;
			16'h3870: y = 16'h200;
			16'h3871: y = 16'h200;
			16'h3872: y = 16'h200;
			16'h3873: y = 16'h200;
			16'h3874: y = 16'h200;
			16'h3875: y = 16'h200;
			16'h3876: y = 16'h200;
			16'h3877: y = 16'h200;
			16'h3878: y = 16'h200;
			16'h3879: y = 16'h200;
			16'h387a: y = 16'h200;
			16'h387b: y = 16'h200;
			16'h387c: y = 16'h200;
			16'h387d: y = 16'h200;
			16'h387e: y = 16'h200;
			16'h387f: y = 16'h200;
			16'h3880: y = 16'h200;
			16'h3881: y = 16'h200;
			16'h3882: y = 16'h200;
			16'h3883: y = 16'h200;
			16'h3884: y = 16'h200;
			16'h3885: y = 16'h200;
			16'h3886: y = 16'h200;
			16'h3887: y = 16'h200;
			16'h3888: y = 16'h200;
			16'h3889: y = 16'h200;
			16'h388a: y = 16'h200;
			16'h388b: y = 16'h200;
			16'h388c: y = 16'h200;
			16'h388d: y = 16'h200;
			16'h388e: y = 16'h200;
			16'h388f: y = 16'h200;
			16'h3890: y = 16'h200;
			16'h3891: y = 16'h200;
			16'h3892: y = 16'h200;
			16'h3893: y = 16'h200;
			16'h3894: y = 16'h200;
			16'h3895: y = 16'h200;
			16'h3896: y = 16'h200;
			16'h3897: y = 16'h200;
			16'h3898: y = 16'h200;
			16'h3899: y = 16'h200;
			16'h389a: y = 16'h200;
			16'h389b: y = 16'h200;
			16'h389c: y = 16'h200;
			16'h389d: y = 16'h200;
			16'h389e: y = 16'h200;
			16'h389f: y = 16'h200;
			16'h38a0: y = 16'h200;
			16'h38a1: y = 16'h200;
			16'h38a2: y = 16'h200;
			16'h38a3: y = 16'h200;
			16'h38a4: y = 16'h200;
			16'h38a5: y = 16'h200;
			16'h38a6: y = 16'h200;
			16'h38a7: y = 16'h200;
			16'h38a8: y = 16'h200;
			16'h38a9: y = 16'h200;
			16'h38aa: y = 16'h200;
			16'h38ab: y = 16'h200;
			16'h38ac: y = 16'h200;
			16'h38ad: y = 16'h200;
			16'h38ae: y = 16'h200;
			16'h38af: y = 16'h200;
			16'h38b0: y = 16'h200;
			16'h38b1: y = 16'h200;
			16'h38b2: y = 16'h200;
			16'h38b3: y = 16'h200;
			16'h38b4: y = 16'h200;
			16'h38b5: y = 16'h200;
			16'h38b6: y = 16'h200;
			16'h38b7: y = 16'h200;
			16'h38b8: y = 16'h200;
			16'h38b9: y = 16'h200;
			16'h38ba: y = 16'h200;
			16'h38bb: y = 16'h200;
			16'h38bc: y = 16'h200;
			16'h38bd: y = 16'h200;
			16'h38be: y = 16'h200;
			16'h38bf: y = 16'h200;
			16'h38c0: y = 16'h200;
			16'h38c1: y = 16'h200;
			16'h38c2: y = 16'h200;
			16'h38c3: y = 16'h200;
			16'h38c4: y = 16'h200;
			16'h38c5: y = 16'h200;
			16'h38c6: y = 16'h200;
			16'h38c7: y = 16'h200;
			16'h38c8: y = 16'h200;
			16'h38c9: y = 16'h200;
			16'h38ca: y = 16'h200;
			16'h38cb: y = 16'h200;
			16'h38cc: y = 16'h200;
			16'h38cd: y = 16'h200;
			16'h38ce: y = 16'h200;
			16'h38cf: y = 16'h200;
			16'h38d0: y = 16'h200;
			16'h38d1: y = 16'h200;
			16'h38d2: y = 16'h200;
			16'h38d3: y = 16'h200;
			16'h38d4: y = 16'h200;
			16'h38d5: y = 16'h200;
			16'h38d6: y = 16'h200;
			16'h38d7: y = 16'h200;
			16'h38d8: y = 16'h200;
			16'h38d9: y = 16'h200;
			16'h38da: y = 16'h200;
			16'h38db: y = 16'h200;
			16'h38dc: y = 16'h200;
			16'h38dd: y = 16'h200;
			16'h38de: y = 16'h200;
			16'h38df: y = 16'h200;
			16'h38e0: y = 16'h200;
			16'h38e1: y = 16'h200;
			16'h38e2: y = 16'h200;
			16'h38e3: y = 16'h200;
			16'h38e4: y = 16'h200;
			16'h38e5: y = 16'h200;
			16'h38e6: y = 16'h200;
			16'h38e7: y = 16'h200;
			16'h38e8: y = 16'h200;
			16'h38e9: y = 16'h200;
			16'h38ea: y = 16'h200;
			16'h38eb: y = 16'h200;
			16'h38ec: y = 16'h200;
			16'h38ed: y = 16'h200;
			16'h38ee: y = 16'h200;
			16'h38ef: y = 16'h200;
			16'h38f0: y = 16'h200;
			16'h38f1: y = 16'h200;
			16'h38f2: y = 16'h200;
			16'h38f3: y = 16'h200;
			16'h38f4: y = 16'h200;
			16'h38f5: y = 16'h200;
			16'h38f6: y = 16'h200;
			16'h38f7: y = 16'h200;
			16'h38f8: y = 16'h200;
			16'h38f9: y = 16'h200;
			16'h38fa: y = 16'h200;
			16'h38fb: y = 16'h200;
			16'h38fc: y = 16'h200;
			16'h38fd: y = 16'h200;
			16'h38fe: y = 16'h200;
			16'h38ff: y = 16'h200;
			16'h3900: y = 16'h200;
			16'h3901: y = 16'h200;
			16'h3902: y = 16'h200;
			16'h3903: y = 16'h200;
			16'h3904: y = 16'h200;
			16'h3905: y = 16'h200;
			16'h3906: y = 16'h200;
			16'h3907: y = 16'h200;
			16'h3908: y = 16'h200;
			16'h3909: y = 16'h200;
			16'h390a: y = 16'h200;
			16'h390b: y = 16'h200;
			16'h390c: y = 16'h200;
			16'h390d: y = 16'h200;
			16'h390e: y = 16'h200;
			16'h390f: y = 16'h200;
			16'h3910: y = 16'h200;
			16'h3911: y = 16'h200;
			16'h3912: y = 16'h200;
			16'h3913: y = 16'h200;
			16'h3914: y = 16'h200;
			16'h3915: y = 16'h200;
			16'h3916: y = 16'h200;
			16'h3917: y = 16'h200;
			16'h3918: y = 16'h200;
			16'h3919: y = 16'h200;
			16'h391a: y = 16'h200;
			16'h391b: y = 16'h200;
			16'h391c: y = 16'h200;
			16'h391d: y = 16'h200;
			16'h391e: y = 16'h200;
			16'h391f: y = 16'h200;
			16'h3920: y = 16'h200;
			16'h3921: y = 16'h200;
			16'h3922: y = 16'h200;
			16'h3923: y = 16'h200;
			16'h3924: y = 16'h200;
			16'h3925: y = 16'h200;
			16'h3926: y = 16'h200;
			16'h3927: y = 16'h200;
			16'h3928: y = 16'h200;
			16'h3929: y = 16'h200;
			16'h392a: y = 16'h200;
			16'h392b: y = 16'h200;
			16'h392c: y = 16'h200;
			16'h392d: y = 16'h200;
			16'h392e: y = 16'h200;
			16'h392f: y = 16'h200;
			16'h3930: y = 16'h200;
			16'h3931: y = 16'h200;
			16'h3932: y = 16'h200;
			16'h3933: y = 16'h200;
			16'h3934: y = 16'h200;
			16'h3935: y = 16'h200;
			16'h3936: y = 16'h200;
			16'h3937: y = 16'h200;
			16'h3938: y = 16'h200;
			16'h3939: y = 16'h200;
			16'h393a: y = 16'h200;
			16'h393b: y = 16'h200;
			16'h393c: y = 16'h200;
			16'h393d: y = 16'h200;
			16'h393e: y = 16'h200;
			16'h393f: y = 16'h200;
			16'h3940: y = 16'h200;
			16'h3941: y = 16'h200;
			16'h3942: y = 16'h200;
			16'h3943: y = 16'h200;
			16'h3944: y = 16'h200;
			16'h3945: y = 16'h200;
			16'h3946: y = 16'h200;
			16'h3947: y = 16'h200;
			16'h3948: y = 16'h200;
			16'h3949: y = 16'h200;
			16'h394a: y = 16'h200;
			16'h394b: y = 16'h200;
			16'h394c: y = 16'h200;
			16'h394d: y = 16'h200;
			16'h394e: y = 16'h200;
			16'h394f: y = 16'h200;
			16'h3950: y = 16'h200;
			16'h3951: y = 16'h200;
			16'h3952: y = 16'h200;
			16'h3953: y = 16'h200;
			16'h3954: y = 16'h200;
			16'h3955: y = 16'h200;
			16'h3956: y = 16'h200;
			16'h3957: y = 16'h200;
			16'h3958: y = 16'h200;
			16'h3959: y = 16'h200;
			16'h395a: y = 16'h200;
			16'h395b: y = 16'h200;
			16'h395c: y = 16'h200;
			16'h395d: y = 16'h200;
			16'h395e: y = 16'h200;
			16'h395f: y = 16'h200;
			16'h3960: y = 16'h200;
			16'h3961: y = 16'h200;
			16'h3962: y = 16'h200;
			16'h3963: y = 16'h200;
			16'h3964: y = 16'h200;
			16'h3965: y = 16'h200;
			16'h3966: y = 16'h200;
			16'h3967: y = 16'h200;
			16'h3968: y = 16'h200;
			16'h3969: y = 16'h200;
			16'h396a: y = 16'h200;
			16'h396b: y = 16'h200;
			16'h396c: y = 16'h200;
			16'h396d: y = 16'h200;
			16'h396e: y = 16'h200;
			16'h396f: y = 16'h200;
			16'h3970: y = 16'h200;
			16'h3971: y = 16'h200;
			16'h3972: y = 16'h200;
			16'h3973: y = 16'h200;
			16'h3974: y = 16'h200;
			16'h3975: y = 16'h200;
			16'h3976: y = 16'h200;
			16'h3977: y = 16'h200;
			16'h3978: y = 16'h200;
			16'h3979: y = 16'h200;
			16'h397a: y = 16'h200;
			16'h397b: y = 16'h200;
			16'h397c: y = 16'h200;
			16'h397d: y = 16'h200;
			16'h397e: y = 16'h200;
			16'h397f: y = 16'h200;
			16'h3980: y = 16'h200;
			16'h3981: y = 16'h200;
			16'h3982: y = 16'h200;
			16'h3983: y = 16'h200;
			16'h3984: y = 16'h200;
			16'h3985: y = 16'h200;
			16'h3986: y = 16'h200;
			16'h3987: y = 16'h200;
			16'h3988: y = 16'h200;
			16'h3989: y = 16'h200;
			16'h398a: y = 16'h200;
			16'h398b: y = 16'h200;
			16'h398c: y = 16'h200;
			16'h398d: y = 16'h200;
			16'h398e: y = 16'h200;
			16'h398f: y = 16'h200;
			16'h3990: y = 16'h200;
			16'h3991: y = 16'h200;
			16'h3992: y = 16'h200;
			16'h3993: y = 16'h200;
			16'h3994: y = 16'h200;
			16'h3995: y = 16'h200;
			16'h3996: y = 16'h200;
			16'h3997: y = 16'h200;
			16'h3998: y = 16'h200;
			16'h3999: y = 16'h200;
			16'h399a: y = 16'h200;
			16'h399b: y = 16'h200;
			16'h399c: y = 16'h200;
			16'h399d: y = 16'h200;
			16'h399e: y = 16'h200;
			16'h399f: y = 16'h200;
			16'h39a0: y = 16'h200;
			16'h39a1: y = 16'h200;
			16'h39a2: y = 16'h200;
			16'h39a3: y = 16'h200;
			16'h39a4: y = 16'h200;
			16'h39a5: y = 16'h200;
			16'h39a6: y = 16'h200;
			16'h39a7: y = 16'h200;
			16'h39a8: y = 16'h200;
			16'h39a9: y = 16'h200;
			16'h39aa: y = 16'h200;
			16'h39ab: y = 16'h200;
			16'h39ac: y = 16'h200;
			16'h39ad: y = 16'h200;
			16'h39ae: y = 16'h200;
			16'h39af: y = 16'h200;
			16'h39b0: y = 16'h200;
			16'h39b1: y = 16'h200;
			16'h39b2: y = 16'h200;
			16'h39b3: y = 16'h200;
			16'h39b4: y = 16'h200;
			16'h39b5: y = 16'h200;
			16'h39b6: y = 16'h200;
			16'h39b7: y = 16'h200;
			16'h39b8: y = 16'h200;
			16'h39b9: y = 16'h200;
			16'h39ba: y = 16'h200;
			16'h39bb: y = 16'h200;
			16'h39bc: y = 16'h200;
			16'h39bd: y = 16'h200;
			16'h39be: y = 16'h200;
			16'h39bf: y = 16'h200;
			16'h39c0: y = 16'h200;
			16'h39c1: y = 16'h200;
			16'h39c2: y = 16'h200;
			16'h39c3: y = 16'h200;
			16'h39c4: y = 16'h200;
			16'h39c5: y = 16'h200;
			16'h39c6: y = 16'h200;
			16'h39c7: y = 16'h200;
			16'h39c8: y = 16'h200;
			16'h39c9: y = 16'h200;
			16'h39ca: y = 16'h200;
			16'h39cb: y = 16'h200;
			16'h39cc: y = 16'h200;
			16'h39cd: y = 16'h200;
			16'h39ce: y = 16'h200;
			16'h39cf: y = 16'h200;
			16'h39d0: y = 16'h200;
			16'h39d1: y = 16'h200;
			16'h39d2: y = 16'h200;
			16'h39d3: y = 16'h200;
			16'h39d4: y = 16'h200;
			16'h39d5: y = 16'h200;
			16'h39d6: y = 16'h200;
			16'h39d7: y = 16'h200;
			16'h39d8: y = 16'h200;
			16'h39d9: y = 16'h200;
			16'h39da: y = 16'h200;
			16'h39db: y = 16'h200;
			16'h39dc: y = 16'h200;
			16'h39dd: y = 16'h200;
			16'h39de: y = 16'h200;
			16'h39df: y = 16'h200;
			16'h39e0: y = 16'h200;
			16'h39e1: y = 16'h200;
			16'h39e2: y = 16'h200;
			16'h39e3: y = 16'h200;
			16'h39e4: y = 16'h200;
			16'h39e5: y = 16'h200;
			16'h39e6: y = 16'h200;
			16'h39e7: y = 16'h200;
			16'h39e8: y = 16'h200;
			16'h39e9: y = 16'h200;
			16'h39ea: y = 16'h200;
			16'h39eb: y = 16'h200;
			16'h39ec: y = 16'h200;
			16'h39ed: y = 16'h200;
			16'h39ee: y = 16'h200;
			16'h39ef: y = 16'h200;
			16'h39f0: y = 16'h200;
			16'h39f1: y = 16'h200;
			16'h39f2: y = 16'h200;
			16'h39f3: y = 16'h200;
			16'h39f4: y = 16'h200;
			16'h39f5: y = 16'h200;
			16'h39f6: y = 16'h200;
			16'h39f7: y = 16'h200;
			16'h39f8: y = 16'h200;
			16'h39f9: y = 16'h200;
			16'h39fa: y = 16'h200;
			16'h39fb: y = 16'h200;
			16'h39fc: y = 16'h200;
			16'h39fd: y = 16'h200;
			16'h39fe: y = 16'h200;
			16'h39ff: y = 16'h200;
			16'h3a00: y = 16'h200;
			16'h3a01: y = 16'h200;
			16'h3a02: y = 16'h200;
			16'h3a03: y = 16'h200;
			16'h3a04: y = 16'h200;
			16'h3a05: y = 16'h200;
			16'h3a06: y = 16'h200;
			16'h3a07: y = 16'h200;
			16'h3a08: y = 16'h200;
			16'h3a09: y = 16'h200;
			16'h3a0a: y = 16'h200;
			16'h3a0b: y = 16'h200;
			16'h3a0c: y = 16'h200;
			16'h3a0d: y = 16'h200;
			16'h3a0e: y = 16'h200;
			16'h3a0f: y = 16'h200;
			16'h3a10: y = 16'h200;
			16'h3a11: y = 16'h200;
			16'h3a12: y = 16'h200;
			16'h3a13: y = 16'h200;
			16'h3a14: y = 16'h200;
			16'h3a15: y = 16'h200;
			16'h3a16: y = 16'h200;
			16'h3a17: y = 16'h200;
			16'h3a18: y = 16'h200;
			16'h3a19: y = 16'h200;
			16'h3a1a: y = 16'h200;
			16'h3a1b: y = 16'h200;
			16'h3a1c: y = 16'h200;
			16'h3a1d: y = 16'h200;
			16'h3a1e: y = 16'h200;
			16'h3a1f: y = 16'h200;
			16'h3a20: y = 16'h200;
			16'h3a21: y = 16'h200;
			16'h3a22: y = 16'h200;
			16'h3a23: y = 16'h200;
			16'h3a24: y = 16'h200;
			16'h3a25: y = 16'h200;
			16'h3a26: y = 16'h200;
			16'h3a27: y = 16'h200;
			16'h3a28: y = 16'h200;
			16'h3a29: y = 16'h200;
			16'h3a2a: y = 16'h200;
			16'h3a2b: y = 16'h200;
			16'h3a2c: y = 16'h200;
			16'h3a2d: y = 16'h200;
			16'h3a2e: y = 16'h200;
			16'h3a2f: y = 16'h200;
			16'h3a30: y = 16'h200;
			16'h3a31: y = 16'h200;
			16'h3a32: y = 16'h200;
			16'h3a33: y = 16'h200;
			16'h3a34: y = 16'h200;
			16'h3a35: y = 16'h200;
			16'h3a36: y = 16'h200;
			16'h3a37: y = 16'h200;
			16'h3a38: y = 16'h200;
			16'h3a39: y = 16'h200;
			16'h3a3a: y = 16'h200;
			16'h3a3b: y = 16'h200;
			16'h3a3c: y = 16'h200;
			16'h3a3d: y = 16'h200;
			16'h3a3e: y = 16'h200;
			16'h3a3f: y = 16'h200;
			16'h3a40: y = 16'h200;
			16'h3a41: y = 16'h200;
			16'h3a42: y = 16'h200;
			16'h3a43: y = 16'h200;
			16'h3a44: y = 16'h200;
			16'h3a45: y = 16'h200;
			16'h3a46: y = 16'h200;
			16'h3a47: y = 16'h200;
			16'h3a48: y = 16'h200;
			16'h3a49: y = 16'h200;
			16'h3a4a: y = 16'h200;
			16'h3a4b: y = 16'h200;
			16'h3a4c: y = 16'h200;
			16'h3a4d: y = 16'h200;
			16'h3a4e: y = 16'h200;
			16'h3a4f: y = 16'h200;
			16'h3a50: y = 16'h200;
			16'h3a51: y = 16'h200;
			16'h3a52: y = 16'h200;
			16'h3a53: y = 16'h200;
			16'h3a54: y = 16'h200;
			16'h3a55: y = 16'h200;
			16'h3a56: y = 16'h200;
			16'h3a57: y = 16'h200;
			16'h3a58: y = 16'h200;
			16'h3a59: y = 16'h200;
			16'h3a5a: y = 16'h200;
			16'h3a5b: y = 16'h200;
			16'h3a5c: y = 16'h200;
			16'h3a5d: y = 16'h200;
			16'h3a5e: y = 16'h200;
			16'h3a5f: y = 16'h200;
			16'h3a60: y = 16'h200;
			16'h3a61: y = 16'h200;
			16'h3a62: y = 16'h200;
			16'h3a63: y = 16'h200;
			16'h3a64: y = 16'h200;
			16'h3a65: y = 16'h200;
			16'h3a66: y = 16'h200;
			16'h3a67: y = 16'h200;
			16'h3a68: y = 16'h200;
			16'h3a69: y = 16'h200;
			16'h3a6a: y = 16'h200;
			16'h3a6b: y = 16'h200;
			16'h3a6c: y = 16'h200;
			16'h3a6d: y = 16'h200;
			16'h3a6e: y = 16'h200;
			16'h3a6f: y = 16'h200;
			16'h3a70: y = 16'h200;
			16'h3a71: y = 16'h200;
			16'h3a72: y = 16'h200;
			16'h3a73: y = 16'h200;
			16'h3a74: y = 16'h200;
			16'h3a75: y = 16'h200;
			16'h3a76: y = 16'h200;
			16'h3a77: y = 16'h200;
			16'h3a78: y = 16'h200;
			16'h3a79: y = 16'h200;
			16'h3a7a: y = 16'h200;
			16'h3a7b: y = 16'h200;
			16'h3a7c: y = 16'h200;
			16'h3a7d: y = 16'h200;
			16'h3a7e: y = 16'h200;
			16'h3a7f: y = 16'h200;
			16'h3a80: y = 16'h200;
			16'h3a81: y = 16'h200;
			16'h3a82: y = 16'h200;
			16'h3a83: y = 16'h200;
			16'h3a84: y = 16'h200;
			16'h3a85: y = 16'h200;
			16'h3a86: y = 16'h200;
			16'h3a87: y = 16'h200;
			16'h3a88: y = 16'h200;
			16'h3a89: y = 16'h200;
			16'h3a8a: y = 16'h200;
			16'h3a8b: y = 16'h200;
			16'h3a8c: y = 16'h200;
			16'h3a8d: y = 16'h200;
			16'h3a8e: y = 16'h200;
			16'h3a8f: y = 16'h200;
			16'h3a90: y = 16'h200;
			16'h3a91: y = 16'h200;
			16'h3a92: y = 16'h200;
			16'h3a93: y = 16'h200;
			16'h3a94: y = 16'h200;
			16'h3a95: y = 16'h200;
			16'h3a96: y = 16'h200;
			16'h3a97: y = 16'h200;
			16'h3a98: y = 16'h200;
			16'h3a99: y = 16'h200;
			16'h3a9a: y = 16'h200;
			16'h3a9b: y = 16'h200;
			16'h3a9c: y = 16'h200;
			16'h3a9d: y = 16'h200;
			16'h3a9e: y = 16'h200;
			16'h3a9f: y = 16'h200;
			16'h3aa0: y = 16'h200;
			16'h3aa1: y = 16'h200;
			16'h3aa2: y = 16'h200;
			16'h3aa3: y = 16'h200;
			16'h3aa4: y = 16'h200;
			16'h3aa5: y = 16'h200;
			16'h3aa6: y = 16'h200;
			16'h3aa7: y = 16'h200;
			16'h3aa8: y = 16'h200;
			16'h3aa9: y = 16'h200;
			16'h3aaa: y = 16'h200;
			16'h3aab: y = 16'h200;
			16'h3aac: y = 16'h200;
			16'h3aad: y = 16'h200;
			16'h3aae: y = 16'h200;
			16'h3aaf: y = 16'h200;
			16'h3ab0: y = 16'h200;
			16'h3ab1: y = 16'h200;
			16'h3ab2: y = 16'h200;
			16'h3ab3: y = 16'h200;
			16'h3ab4: y = 16'h200;
			16'h3ab5: y = 16'h200;
			16'h3ab6: y = 16'h200;
			16'h3ab7: y = 16'h200;
			16'h3ab8: y = 16'h200;
			16'h3ab9: y = 16'h200;
			16'h3aba: y = 16'h200;
			16'h3abb: y = 16'h200;
			16'h3abc: y = 16'h200;
			16'h3abd: y = 16'h200;
			16'h3abe: y = 16'h200;
			16'h3abf: y = 16'h200;
			16'h3ac0: y = 16'h200;
			16'h3ac1: y = 16'h200;
			16'h3ac2: y = 16'h200;
			16'h3ac3: y = 16'h200;
			16'h3ac4: y = 16'h200;
			16'h3ac5: y = 16'h200;
			16'h3ac6: y = 16'h200;
			16'h3ac7: y = 16'h200;
			16'h3ac8: y = 16'h200;
			16'h3ac9: y = 16'h200;
			16'h3aca: y = 16'h200;
			16'h3acb: y = 16'h200;
			16'h3acc: y = 16'h200;
			16'h3acd: y = 16'h200;
			16'h3ace: y = 16'h200;
			16'h3acf: y = 16'h200;
			16'h3ad0: y = 16'h200;
			16'h3ad1: y = 16'h200;
			16'h3ad2: y = 16'h200;
			16'h3ad3: y = 16'h200;
			16'h3ad4: y = 16'h200;
			16'h3ad5: y = 16'h200;
			16'h3ad6: y = 16'h200;
			16'h3ad7: y = 16'h200;
			16'h3ad8: y = 16'h200;
			16'h3ad9: y = 16'h200;
			16'h3ada: y = 16'h200;
			16'h3adb: y = 16'h200;
			16'h3adc: y = 16'h200;
			16'h3add: y = 16'h200;
			16'h3ade: y = 16'h200;
			16'h3adf: y = 16'h200;
			16'h3ae0: y = 16'h200;
			16'h3ae1: y = 16'h200;
			16'h3ae2: y = 16'h200;
			16'h3ae3: y = 16'h200;
			16'h3ae4: y = 16'h200;
			16'h3ae5: y = 16'h200;
			16'h3ae6: y = 16'h200;
			16'h3ae7: y = 16'h200;
			16'h3ae8: y = 16'h200;
			16'h3ae9: y = 16'h200;
			16'h3aea: y = 16'h200;
			16'h3aeb: y = 16'h200;
			16'h3aec: y = 16'h200;
			16'h3aed: y = 16'h200;
			16'h3aee: y = 16'h200;
			16'h3aef: y = 16'h200;
			16'h3af0: y = 16'h200;
			16'h3af1: y = 16'h200;
			16'h3af2: y = 16'h200;
			16'h3af3: y = 16'h200;
			16'h3af4: y = 16'h200;
			16'h3af5: y = 16'h200;
			16'h3af6: y = 16'h200;
			16'h3af7: y = 16'h200;
			16'h3af8: y = 16'h200;
			16'h3af9: y = 16'h200;
			16'h3afa: y = 16'h200;
			16'h3afb: y = 16'h200;
			16'h3afc: y = 16'h200;
			16'h3afd: y = 16'h200;
			16'h3afe: y = 16'h200;
			16'h3aff: y = 16'h200;
			16'h3b00: y = 16'h200;
			16'h3b01: y = 16'h200;
			16'h3b02: y = 16'h200;
			16'h3b03: y = 16'h200;
			16'h3b04: y = 16'h200;
			16'h3b05: y = 16'h200;
			16'h3b06: y = 16'h200;
			16'h3b07: y = 16'h200;
			16'h3b08: y = 16'h200;
			16'h3b09: y = 16'h200;
			16'h3b0a: y = 16'h200;
			16'h3b0b: y = 16'h200;
			16'h3b0c: y = 16'h200;
			16'h3b0d: y = 16'h200;
			16'h3b0e: y = 16'h200;
			16'h3b0f: y = 16'h200;
			16'h3b10: y = 16'h200;
			16'h3b11: y = 16'h200;
			16'h3b12: y = 16'h200;
			16'h3b13: y = 16'h200;
			16'h3b14: y = 16'h200;
			16'h3b15: y = 16'h200;
			16'h3b16: y = 16'h200;
			16'h3b17: y = 16'h200;
			16'h3b18: y = 16'h200;
			16'h3b19: y = 16'h200;
			16'h3b1a: y = 16'h200;
			16'h3b1b: y = 16'h200;
			16'h3b1c: y = 16'h200;
			16'h3b1d: y = 16'h200;
			16'h3b1e: y = 16'h200;
			16'h3b1f: y = 16'h200;
			16'h3b20: y = 16'h200;
			16'h3b21: y = 16'h200;
			16'h3b22: y = 16'h200;
			16'h3b23: y = 16'h200;
			16'h3b24: y = 16'h200;
			16'h3b25: y = 16'h200;
			16'h3b26: y = 16'h200;
			16'h3b27: y = 16'h200;
			16'h3b28: y = 16'h200;
			16'h3b29: y = 16'h200;
			16'h3b2a: y = 16'h200;
			16'h3b2b: y = 16'h200;
			16'h3b2c: y = 16'h200;
			16'h3b2d: y = 16'h200;
			16'h3b2e: y = 16'h200;
			16'h3b2f: y = 16'h200;
			16'h3b30: y = 16'h200;
			16'h3b31: y = 16'h200;
			16'h3b32: y = 16'h200;
			16'h3b33: y = 16'h200;
			16'h3b34: y = 16'h200;
			16'h3b35: y = 16'h200;
			16'h3b36: y = 16'h200;
			16'h3b37: y = 16'h200;
			16'h3b38: y = 16'h200;
			16'h3b39: y = 16'h200;
			16'h3b3a: y = 16'h200;
			16'h3b3b: y = 16'h200;
			16'h3b3c: y = 16'h200;
			16'h3b3d: y = 16'h200;
			16'h3b3e: y = 16'h200;
			16'h3b3f: y = 16'h200;
			16'h3b40: y = 16'h200;
			16'h3b41: y = 16'h200;
			16'h3b42: y = 16'h200;
			16'h3b43: y = 16'h200;
			16'h3b44: y = 16'h200;
			16'h3b45: y = 16'h200;
			16'h3b46: y = 16'h200;
			16'h3b47: y = 16'h200;
			16'h3b48: y = 16'h200;
			16'h3b49: y = 16'h200;
			16'h3b4a: y = 16'h200;
			16'h3b4b: y = 16'h200;
			16'h3b4c: y = 16'h200;
			16'h3b4d: y = 16'h200;
			16'h3b4e: y = 16'h200;
			16'h3b4f: y = 16'h200;
			16'h3b50: y = 16'h200;
			16'h3b51: y = 16'h200;
			16'h3b52: y = 16'h200;
			16'h3b53: y = 16'h200;
			16'h3b54: y = 16'h200;
			16'h3b55: y = 16'h200;
			16'h3b56: y = 16'h200;
			16'h3b57: y = 16'h200;
			16'h3b58: y = 16'h200;
			16'h3b59: y = 16'h200;
			16'h3b5a: y = 16'h200;
			16'h3b5b: y = 16'h200;
			16'h3b5c: y = 16'h200;
			16'h3b5d: y = 16'h200;
			16'h3b5e: y = 16'h200;
			16'h3b5f: y = 16'h200;
			16'h3b60: y = 16'h200;
			16'h3b61: y = 16'h200;
			16'h3b62: y = 16'h200;
			16'h3b63: y = 16'h200;
			16'h3b64: y = 16'h200;
			16'h3b65: y = 16'h200;
			16'h3b66: y = 16'h200;
			16'h3b67: y = 16'h200;
			16'h3b68: y = 16'h200;
			16'h3b69: y = 16'h200;
			16'h3b6a: y = 16'h200;
			16'h3b6b: y = 16'h200;
			16'h3b6c: y = 16'h200;
			16'h3b6d: y = 16'h200;
			16'h3b6e: y = 16'h200;
			16'h3b6f: y = 16'h200;
			16'h3b70: y = 16'h200;
			16'h3b71: y = 16'h200;
			16'h3b72: y = 16'h200;
			16'h3b73: y = 16'h200;
			16'h3b74: y = 16'h200;
			16'h3b75: y = 16'h200;
			16'h3b76: y = 16'h200;
			16'h3b77: y = 16'h200;
			16'h3b78: y = 16'h200;
			16'h3b79: y = 16'h200;
			16'h3b7a: y = 16'h200;
			16'h3b7b: y = 16'h200;
			16'h3b7c: y = 16'h200;
			16'h3b7d: y = 16'h200;
			16'h3b7e: y = 16'h200;
			16'h3b7f: y = 16'h200;
			16'h3b80: y = 16'h200;
			16'h3b81: y = 16'h200;
			16'h3b82: y = 16'h200;
			16'h3b83: y = 16'h200;
			16'h3b84: y = 16'h200;
			16'h3b85: y = 16'h200;
			16'h3b86: y = 16'h200;
			16'h3b87: y = 16'h200;
			16'h3b88: y = 16'h200;
			16'h3b89: y = 16'h200;
			16'h3b8a: y = 16'h200;
			16'h3b8b: y = 16'h200;
			16'h3b8c: y = 16'h200;
			16'h3b8d: y = 16'h200;
			16'h3b8e: y = 16'h200;
			16'h3b8f: y = 16'h200;
			16'h3b90: y = 16'h200;
			16'h3b91: y = 16'h200;
			16'h3b92: y = 16'h200;
			16'h3b93: y = 16'h200;
			16'h3b94: y = 16'h200;
			16'h3b95: y = 16'h200;
			16'h3b96: y = 16'h200;
			16'h3b97: y = 16'h200;
			16'h3b98: y = 16'h200;
			16'h3b99: y = 16'h200;
			16'h3b9a: y = 16'h200;
			16'h3b9b: y = 16'h200;
			16'h3b9c: y = 16'h200;
			16'h3b9d: y = 16'h200;
			16'h3b9e: y = 16'h200;
			16'h3b9f: y = 16'h200;
			16'h3ba0: y = 16'h200;
			16'h3ba1: y = 16'h200;
			16'h3ba2: y = 16'h200;
			16'h3ba3: y = 16'h200;
			16'h3ba4: y = 16'h200;
			16'h3ba5: y = 16'h200;
			16'h3ba6: y = 16'h200;
			16'h3ba7: y = 16'h200;
			16'h3ba8: y = 16'h200;
			16'h3ba9: y = 16'h200;
			16'h3baa: y = 16'h200;
			16'h3bab: y = 16'h200;
			16'h3bac: y = 16'h200;
			16'h3bad: y = 16'h200;
			16'h3bae: y = 16'h200;
			16'h3baf: y = 16'h200;
			16'h3bb0: y = 16'h200;
			16'h3bb1: y = 16'h200;
			16'h3bb2: y = 16'h200;
			16'h3bb3: y = 16'h200;
			16'h3bb4: y = 16'h200;
			16'h3bb5: y = 16'h200;
			16'h3bb6: y = 16'h200;
			16'h3bb7: y = 16'h200;
			16'h3bb8: y = 16'h200;
			16'h3bb9: y = 16'h200;
			16'h3bba: y = 16'h200;
			16'h3bbb: y = 16'h200;
			16'h3bbc: y = 16'h200;
			16'h3bbd: y = 16'h200;
			16'h3bbe: y = 16'h200;
			16'h3bbf: y = 16'h200;
			16'h3bc0: y = 16'h200;
			16'h3bc1: y = 16'h200;
			16'h3bc2: y = 16'h200;
			16'h3bc3: y = 16'h200;
			16'h3bc4: y = 16'h200;
			16'h3bc5: y = 16'h200;
			16'h3bc6: y = 16'h200;
			16'h3bc7: y = 16'h200;
			16'h3bc8: y = 16'h200;
			16'h3bc9: y = 16'h200;
			16'h3bca: y = 16'h200;
			16'h3bcb: y = 16'h200;
			16'h3bcc: y = 16'h200;
			16'h3bcd: y = 16'h200;
			16'h3bce: y = 16'h200;
			16'h3bcf: y = 16'h200;
			16'h3bd0: y = 16'h200;
			16'h3bd1: y = 16'h200;
			16'h3bd2: y = 16'h200;
			16'h3bd3: y = 16'h200;
			16'h3bd4: y = 16'h200;
			16'h3bd5: y = 16'h200;
			16'h3bd6: y = 16'h200;
			16'h3bd7: y = 16'h200;
			16'h3bd8: y = 16'h200;
			16'h3bd9: y = 16'h200;
			16'h3bda: y = 16'h200;
			16'h3bdb: y = 16'h200;
			16'h3bdc: y = 16'h200;
			16'h3bdd: y = 16'h200;
			16'h3bde: y = 16'h200;
			16'h3bdf: y = 16'h200;
			16'h3be0: y = 16'h200;
			16'h3be1: y = 16'h200;
			16'h3be2: y = 16'h200;
			16'h3be3: y = 16'h200;
			16'h3be4: y = 16'h200;
			16'h3be5: y = 16'h200;
			16'h3be6: y = 16'h200;
			16'h3be7: y = 16'h200;
			16'h3be8: y = 16'h200;
			16'h3be9: y = 16'h200;
			16'h3bea: y = 16'h200;
			16'h3beb: y = 16'h200;
			16'h3bec: y = 16'h200;
			16'h3bed: y = 16'h200;
			16'h3bee: y = 16'h200;
			16'h3bef: y = 16'h200;
			16'h3bf0: y = 16'h200;
			16'h3bf1: y = 16'h200;
			16'h3bf2: y = 16'h200;
			16'h3bf3: y = 16'h200;
			16'h3bf4: y = 16'h200;
			16'h3bf5: y = 16'h200;
			16'h3bf6: y = 16'h200;
			16'h3bf7: y = 16'h200;
			16'h3bf8: y = 16'h200;
			16'h3bf9: y = 16'h200;
			16'h3bfa: y = 16'h200;
			16'h3bfb: y = 16'h200;
			16'h3bfc: y = 16'h200;
			16'h3bfd: y = 16'h200;
			16'h3bfe: y = 16'h200;
			16'h3bff: y = 16'h200;
			16'h3c00: y = 16'h200;
			16'h3c01: y = 16'h200;
			16'h3c02: y = 16'h200;
			16'h3c03: y = 16'h200;
			16'h3c04: y = 16'h200;
			16'h3c05: y = 16'h200;
			16'h3c06: y = 16'h200;
			16'h3c07: y = 16'h200;
			16'h3c08: y = 16'h200;
			16'h3c09: y = 16'h200;
			16'h3c0a: y = 16'h200;
			16'h3c0b: y = 16'h200;
			16'h3c0c: y = 16'h200;
			16'h3c0d: y = 16'h200;
			16'h3c0e: y = 16'h200;
			16'h3c0f: y = 16'h200;
			16'h3c10: y = 16'h200;
			16'h3c11: y = 16'h200;
			16'h3c12: y = 16'h200;
			16'h3c13: y = 16'h200;
			16'h3c14: y = 16'h200;
			16'h3c15: y = 16'h200;
			16'h3c16: y = 16'h200;
			16'h3c17: y = 16'h200;
			16'h3c18: y = 16'h200;
			16'h3c19: y = 16'h200;
			16'h3c1a: y = 16'h200;
			16'h3c1b: y = 16'h200;
			16'h3c1c: y = 16'h200;
			16'h3c1d: y = 16'h200;
			16'h3c1e: y = 16'h200;
			16'h3c1f: y = 16'h200;
			16'h3c20: y = 16'h200;
			16'h3c21: y = 16'h200;
			16'h3c22: y = 16'h200;
			16'h3c23: y = 16'h200;
			16'h3c24: y = 16'h200;
			16'h3c25: y = 16'h200;
			16'h3c26: y = 16'h200;
			16'h3c27: y = 16'h200;
			16'h3c28: y = 16'h200;
			16'h3c29: y = 16'h200;
			16'h3c2a: y = 16'h200;
			16'h3c2b: y = 16'h200;
			16'h3c2c: y = 16'h200;
			16'h3c2d: y = 16'h200;
			16'h3c2e: y = 16'h200;
			16'h3c2f: y = 16'h200;
			16'h3c30: y = 16'h200;
			16'h3c31: y = 16'h200;
			16'h3c32: y = 16'h200;
			16'h3c33: y = 16'h200;
			16'h3c34: y = 16'h200;
			16'h3c35: y = 16'h200;
			16'h3c36: y = 16'h200;
			16'h3c37: y = 16'h200;
			16'h3c38: y = 16'h200;
			16'h3c39: y = 16'h200;
			16'h3c3a: y = 16'h200;
			16'h3c3b: y = 16'h200;
			16'h3c3c: y = 16'h200;
			16'h3c3d: y = 16'h200;
			16'h3c3e: y = 16'h200;
			16'h3c3f: y = 16'h200;
			16'h3c40: y = 16'h200;
			16'h3c41: y = 16'h200;
			16'h3c42: y = 16'h200;
			16'h3c43: y = 16'h200;
			16'h3c44: y = 16'h200;
			16'h3c45: y = 16'h200;
			16'h3c46: y = 16'h200;
			16'h3c47: y = 16'h200;
			16'h3c48: y = 16'h200;
			16'h3c49: y = 16'h200;
			16'h3c4a: y = 16'h200;
			16'h3c4b: y = 16'h200;
			16'h3c4c: y = 16'h200;
			16'h3c4d: y = 16'h200;
			16'h3c4e: y = 16'h200;
			16'h3c4f: y = 16'h200;
			16'h3c50: y = 16'h200;
			16'h3c51: y = 16'h200;
			16'h3c52: y = 16'h200;
			16'h3c53: y = 16'h200;
			16'h3c54: y = 16'h200;
			16'h3c55: y = 16'h200;
			16'h3c56: y = 16'h200;
			16'h3c57: y = 16'h200;
			16'h3c58: y = 16'h200;
			16'h3c59: y = 16'h200;
			16'h3c5a: y = 16'h200;
			16'h3c5b: y = 16'h200;
			16'h3c5c: y = 16'h200;
			16'h3c5d: y = 16'h200;
			16'h3c5e: y = 16'h200;
			16'h3c5f: y = 16'h200;
			16'h3c60: y = 16'h200;
			16'h3c61: y = 16'h200;
			16'h3c62: y = 16'h200;
			16'h3c63: y = 16'h200;
			16'h3c64: y = 16'h200;
			16'h3c65: y = 16'h200;
			16'h3c66: y = 16'h200;
			16'h3c67: y = 16'h200;
			16'h3c68: y = 16'h200;
			16'h3c69: y = 16'h200;
			16'h3c6a: y = 16'h200;
			16'h3c6b: y = 16'h200;
			16'h3c6c: y = 16'h200;
			16'h3c6d: y = 16'h200;
			16'h3c6e: y = 16'h200;
			16'h3c6f: y = 16'h200;
			16'h3c70: y = 16'h200;
			16'h3c71: y = 16'h200;
			16'h3c72: y = 16'h200;
			16'h3c73: y = 16'h200;
			16'h3c74: y = 16'h200;
			16'h3c75: y = 16'h200;
			16'h3c76: y = 16'h200;
			16'h3c77: y = 16'h200;
			16'h3c78: y = 16'h200;
			16'h3c79: y = 16'h200;
			16'h3c7a: y = 16'h200;
			16'h3c7b: y = 16'h200;
			16'h3c7c: y = 16'h200;
			16'h3c7d: y = 16'h200;
			16'h3c7e: y = 16'h200;
			16'h3c7f: y = 16'h200;
			16'h3c80: y = 16'h200;
			16'h3c81: y = 16'h200;
			16'h3c82: y = 16'h200;
			16'h3c83: y = 16'h200;
			16'h3c84: y = 16'h200;
			16'h3c85: y = 16'h200;
			16'h3c86: y = 16'h200;
			16'h3c87: y = 16'h200;
			16'h3c88: y = 16'h200;
			16'h3c89: y = 16'h200;
			16'h3c8a: y = 16'h200;
			16'h3c8b: y = 16'h200;
			16'h3c8c: y = 16'h200;
			16'h3c8d: y = 16'h200;
			16'h3c8e: y = 16'h200;
			16'h3c8f: y = 16'h200;
			16'h3c90: y = 16'h200;
			16'h3c91: y = 16'h200;
			16'h3c92: y = 16'h200;
			16'h3c93: y = 16'h200;
			16'h3c94: y = 16'h200;
			16'h3c95: y = 16'h200;
			16'h3c96: y = 16'h200;
			16'h3c97: y = 16'h200;
			16'h3c98: y = 16'h200;
			16'h3c99: y = 16'h200;
			16'h3c9a: y = 16'h200;
			16'h3c9b: y = 16'h200;
			16'h3c9c: y = 16'h200;
			16'h3c9d: y = 16'h200;
			16'h3c9e: y = 16'h200;
			16'h3c9f: y = 16'h200;
			16'h3ca0: y = 16'h200;
			16'h3ca1: y = 16'h200;
			16'h3ca2: y = 16'h200;
			16'h3ca3: y = 16'h200;
			16'h3ca4: y = 16'h200;
			16'h3ca5: y = 16'h200;
			16'h3ca6: y = 16'h200;
			16'h3ca7: y = 16'h200;
			16'h3ca8: y = 16'h200;
			16'h3ca9: y = 16'h200;
			16'h3caa: y = 16'h200;
			16'h3cab: y = 16'h200;
			16'h3cac: y = 16'h200;
			16'h3cad: y = 16'h200;
			16'h3cae: y = 16'h200;
			16'h3caf: y = 16'h200;
			16'h3cb0: y = 16'h200;
			16'h3cb1: y = 16'h200;
			16'h3cb2: y = 16'h200;
			16'h3cb3: y = 16'h200;
			16'h3cb4: y = 16'h200;
			16'h3cb5: y = 16'h200;
			16'h3cb6: y = 16'h200;
			16'h3cb7: y = 16'h200;
			16'h3cb8: y = 16'h200;
			16'h3cb9: y = 16'h200;
			16'h3cba: y = 16'h200;
			16'h3cbb: y = 16'h200;
			16'h3cbc: y = 16'h200;
			16'h3cbd: y = 16'h200;
			16'h3cbe: y = 16'h200;
			16'h3cbf: y = 16'h200;
			16'h3cc0: y = 16'h200;
			16'h3cc1: y = 16'h200;
			16'h3cc2: y = 16'h200;
			16'h3cc3: y = 16'h200;
			16'h3cc4: y = 16'h200;
			16'h3cc5: y = 16'h200;
			16'h3cc6: y = 16'h200;
			16'h3cc7: y = 16'h200;
			16'h3cc8: y = 16'h200;
			16'h3cc9: y = 16'h200;
			16'h3cca: y = 16'h200;
			16'h3ccb: y = 16'h200;
			16'h3ccc: y = 16'h200;
			16'h3ccd: y = 16'h200;
			16'h3cce: y = 16'h200;
			16'h3ccf: y = 16'h200;
			16'h3cd0: y = 16'h200;
			16'h3cd1: y = 16'h200;
			16'h3cd2: y = 16'h200;
			16'h3cd3: y = 16'h200;
			16'h3cd4: y = 16'h200;
			16'h3cd5: y = 16'h200;
			16'h3cd6: y = 16'h200;
			16'h3cd7: y = 16'h200;
			16'h3cd8: y = 16'h200;
			16'h3cd9: y = 16'h200;
			16'h3cda: y = 16'h200;
			16'h3cdb: y = 16'h200;
			16'h3cdc: y = 16'h200;
			16'h3cdd: y = 16'h200;
			16'h3cde: y = 16'h200;
			16'h3cdf: y = 16'h200;
			16'h3ce0: y = 16'h200;
			16'h3ce1: y = 16'h200;
			16'h3ce2: y = 16'h200;
			16'h3ce3: y = 16'h200;
			16'h3ce4: y = 16'h200;
			16'h3ce5: y = 16'h200;
			16'h3ce6: y = 16'h200;
			16'h3ce7: y = 16'h200;
			16'h3ce8: y = 16'h200;
			16'h3ce9: y = 16'h200;
			16'h3cea: y = 16'h200;
			16'h3ceb: y = 16'h200;
			16'h3cec: y = 16'h200;
			16'h3ced: y = 16'h200;
			16'h3cee: y = 16'h200;
			16'h3cef: y = 16'h200;
			16'h3cf0: y = 16'h200;
			16'h3cf1: y = 16'h200;
			16'h3cf2: y = 16'h200;
			16'h3cf3: y = 16'h200;
			16'h3cf4: y = 16'h200;
			16'h3cf5: y = 16'h200;
			16'h3cf6: y = 16'h200;
			16'h3cf7: y = 16'h200;
			16'h3cf8: y = 16'h200;
			16'h3cf9: y = 16'h200;
			16'h3cfa: y = 16'h200;
			16'h3cfb: y = 16'h200;
			16'h3cfc: y = 16'h200;
			16'h3cfd: y = 16'h200;
			16'h3cfe: y = 16'h200;
			16'h3cff: y = 16'h200;
			16'h3d00: y = 16'h200;
			16'h3d01: y = 16'h200;
			16'h3d02: y = 16'h200;
			16'h3d03: y = 16'h200;
			16'h3d04: y = 16'h200;
			16'h3d05: y = 16'h200;
			16'h3d06: y = 16'h200;
			16'h3d07: y = 16'h200;
			16'h3d08: y = 16'h200;
			16'h3d09: y = 16'h200;
			16'h3d0a: y = 16'h200;
			16'h3d0b: y = 16'h200;
			16'h3d0c: y = 16'h200;
			16'h3d0d: y = 16'h200;
			16'h3d0e: y = 16'h200;
			16'h3d0f: y = 16'h200;
			16'h3d10: y = 16'h200;
			16'h3d11: y = 16'h200;
			16'h3d12: y = 16'h200;
			16'h3d13: y = 16'h200;
			16'h3d14: y = 16'h200;
			16'h3d15: y = 16'h200;
			16'h3d16: y = 16'h200;
			16'h3d17: y = 16'h200;
			16'h3d18: y = 16'h200;
			16'h3d19: y = 16'h200;
			16'h3d1a: y = 16'h200;
			16'h3d1b: y = 16'h200;
			16'h3d1c: y = 16'h200;
			16'h3d1d: y = 16'h200;
			16'h3d1e: y = 16'h200;
			16'h3d1f: y = 16'h200;
			16'h3d20: y = 16'h200;
			16'h3d21: y = 16'h200;
			16'h3d22: y = 16'h200;
			16'h3d23: y = 16'h200;
			16'h3d24: y = 16'h200;
			16'h3d25: y = 16'h200;
			16'h3d26: y = 16'h200;
			16'h3d27: y = 16'h200;
			16'h3d28: y = 16'h200;
			16'h3d29: y = 16'h200;
			16'h3d2a: y = 16'h200;
			16'h3d2b: y = 16'h200;
			16'h3d2c: y = 16'h200;
			16'h3d2d: y = 16'h200;
			16'h3d2e: y = 16'h200;
			16'h3d2f: y = 16'h200;
			16'h3d30: y = 16'h200;
			16'h3d31: y = 16'h200;
			16'h3d32: y = 16'h200;
			16'h3d33: y = 16'h200;
			16'h3d34: y = 16'h200;
			16'h3d35: y = 16'h200;
			16'h3d36: y = 16'h200;
			16'h3d37: y = 16'h200;
			16'h3d38: y = 16'h200;
			16'h3d39: y = 16'h200;
			16'h3d3a: y = 16'h200;
			16'h3d3b: y = 16'h200;
			16'h3d3c: y = 16'h200;
			16'h3d3d: y = 16'h200;
			16'h3d3e: y = 16'h200;
			16'h3d3f: y = 16'h200;
			16'h3d40: y = 16'h200;
			16'h3d41: y = 16'h200;
			16'h3d42: y = 16'h200;
			16'h3d43: y = 16'h200;
			16'h3d44: y = 16'h200;
			16'h3d45: y = 16'h200;
			16'h3d46: y = 16'h200;
			16'h3d47: y = 16'h200;
			16'h3d48: y = 16'h200;
			16'h3d49: y = 16'h200;
			16'h3d4a: y = 16'h200;
			16'h3d4b: y = 16'h200;
			16'h3d4c: y = 16'h200;
			16'h3d4d: y = 16'h200;
			16'h3d4e: y = 16'h200;
			16'h3d4f: y = 16'h200;
			16'h3d50: y = 16'h200;
			16'h3d51: y = 16'h200;
			16'h3d52: y = 16'h200;
			16'h3d53: y = 16'h200;
			16'h3d54: y = 16'h200;
			16'h3d55: y = 16'h200;
			16'h3d56: y = 16'h200;
			16'h3d57: y = 16'h200;
			16'h3d58: y = 16'h200;
			16'h3d59: y = 16'h200;
			16'h3d5a: y = 16'h200;
			16'h3d5b: y = 16'h200;
			16'h3d5c: y = 16'h200;
			16'h3d5d: y = 16'h200;
			16'h3d5e: y = 16'h200;
			16'h3d5f: y = 16'h200;
			16'h3d60: y = 16'h200;
			16'h3d61: y = 16'h200;
			16'h3d62: y = 16'h200;
			16'h3d63: y = 16'h200;
			16'h3d64: y = 16'h200;
			16'h3d65: y = 16'h200;
			16'h3d66: y = 16'h200;
			16'h3d67: y = 16'h200;
			16'h3d68: y = 16'h200;
			16'h3d69: y = 16'h200;
			16'h3d6a: y = 16'h200;
			16'h3d6b: y = 16'h200;
			16'h3d6c: y = 16'h200;
			16'h3d6d: y = 16'h200;
			16'h3d6e: y = 16'h200;
			16'h3d6f: y = 16'h200;
			16'h3d70: y = 16'h200;
			16'h3d71: y = 16'h200;
			16'h3d72: y = 16'h200;
			16'h3d73: y = 16'h200;
			16'h3d74: y = 16'h200;
			16'h3d75: y = 16'h200;
			16'h3d76: y = 16'h200;
			16'h3d77: y = 16'h200;
			16'h3d78: y = 16'h200;
			16'h3d79: y = 16'h200;
			16'h3d7a: y = 16'h200;
			16'h3d7b: y = 16'h200;
			16'h3d7c: y = 16'h200;
			16'h3d7d: y = 16'h200;
			16'h3d7e: y = 16'h200;
			16'h3d7f: y = 16'h200;
			16'h3d80: y = 16'h200;
			16'h3d81: y = 16'h200;
			16'h3d82: y = 16'h200;
			16'h3d83: y = 16'h200;
			16'h3d84: y = 16'h200;
			16'h3d85: y = 16'h200;
			16'h3d86: y = 16'h200;
			16'h3d87: y = 16'h200;
			16'h3d88: y = 16'h200;
			16'h3d89: y = 16'h200;
			16'h3d8a: y = 16'h200;
			16'h3d8b: y = 16'h200;
			16'h3d8c: y = 16'h200;
			16'h3d8d: y = 16'h200;
			16'h3d8e: y = 16'h200;
			16'h3d8f: y = 16'h200;
			16'h3d90: y = 16'h200;
			16'h3d91: y = 16'h200;
			16'h3d92: y = 16'h200;
			16'h3d93: y = 16'h200;
			16'h3d94: y = 16'h200;
			16'h3d95: y = 16'h200;
			16'h3d96: y = 16'h200;
			16'h3d97: y = 16'h200;
			16'h3d98: y = 16'h200;
			16'h3d99: y = 16'h200;
			16'h3d9a: y = 16'h200;
			16'h3d9b: y = 16'h200;
			16'h3d9c: y = 16'h200;
			16'h3d9d: y = 16'h200;
			16'h3d9e: y = 16'h200;
			16'h3d9f: y = 16'h200;
			16'h3da0: y = 16'h200;
			16'h3da1: y = 16'h200;
			16'h3da2: y = 16'h200;
			16'h3da3: y = 16'h200;
			16'h3da4: y = 16'h200;
			16'h3da5: y = 16'h200;
			16'h3da6: y = 16'h200;
			16'h3da7: y = 16'h200;
			16'h3da8: y = 16'h200;
			16'h3da9: y = 16'h200;
			16'h3daa: y = 16'h200;
			16'h3dab: y = 16'h200;
			16'h3dac: y = 16'h200;
			16'h3dad: y = 16'h200;
			16'h3dae: y = 16'h200;
			16'h3daf: y = 16'h200;
			16'h3db0: y = 16'h200;
			16'h3db1: y = 16'h200;
			16'h3db2: y = 16'h200;
			16'h3db3: y = 16'h200;
			16'h3db4: y = 16'h200;
			16'h3db5: y = 16'h200;
			16'h3db6: y = 16'h200;
			16'h3db7: y = 16'h200;
			16'h3db8: y = 16'h200;
			16'h3db9: y = 16'h200;
			16'h3dba: y = 16'h200;
			16'h3dbb: y = 16'h200;
			16'h3dbc: y = 16'h200;
			16'h3dbd: y = 16'h200;
			16'h3dbe: y = 16'h200;
			16'h3dbf: y = 16'h200;
			16'h3dc0: y = 16'h200;
			16'h3dc1: y = 16'h200;
			16'h3dc2: y = 16'h200;
			16'h3dc3: y = 16'h200;
			16'h3dc4: y = 16'h200;
			16'h3dc5: y = 16'h200;
			16'h3dc6: y = 16'h200;
			16'h3dc7: y = 16'h200;
			16'h3dc8: y = 16'h200;
			16'h3dc9: y = 16'h200;
			16'h3dca: y = 16'h200;
			16'h3dcb: y = 16'h200;
			16'h3dcc: y = 16'h200;
			16'h3dcd: y = 16'h200;
			16'h3dce: y = 16'h200;
			16'h3dcf: y = 16'h200;
			16'h3dd0: y = 16'h200;
			16'h3dd1: y = 16'h200;
			16'h3dd2: y = 16'h200;
			16'h3dd3: y = 16'h200;
			16'h3dd4: y = 16'h200;
			16'h3dd5: y = 16'h200;
			16'h3dd6: y = 16'h200;
			16'h3dd7: y = 16'h200;
			16'h3dd8: y = 16'h200;
			16'h3dd9: y = 16'h200;
			16'h3dda: y = 16'h200;
			16'h3ddb: y = 16'h200;
			16'h3ddc: y = 16'h200;
			16'h3ddd: y = 16'h200;
			16'h3dde: y = 16'h200;
			16'h3ddf: y = 16'h200;
			16'h3de0: y = 16'h200;
			16'h3de1: y = 16'h200;
			16'h3de2: y = 16'h200;
			16'h3de3: y = 16'h200;
			16'h3de4: y = 16'h200;
			16'h3de5: y = 16'h200;
			16'h3de6: y = 16'h200;
			16'h3de7: y = 16'h200;
			16'h3de8: y = 16'h200;
			16'h3de9: y = 16'h200;
			16'h3dea: y = 16'h200;
			16'h3deb: y = 16'h200;
			16'h3dec: y = 16'h200;
			16'h3ded: y = 16'h200;
			16'h3dee: y = 16'h200;
			16'h3def: y = 16'h200;
			16'h3df0: y = 16'h200;
			16'h3df1: y = 16'h200;
			16'h3df2: y = 16'h200;
			16'h3df3: y = 16'h200;
			16'h3df4: y = 16'h200;
			16'h3df5: y = 16'h200;
			16'h3df6: y = 16'h200;
			16'h3df7: y = 16'h200;
			16'h3df8: y = 16'h200;
			16'h3df9: y = 16'h200;
			16'h3dfa: y = 16'h200;
			16'h3dfb: y = 16'h200;
			16'h3dfc: y = 16'h200;
			16'h3dfd: y = 16'h200;
			16'h3dfe: y = 16'h200;
			16'h3dff: y = 16'h200;
			16'h3e00: y = 16'h200;
			16'h3e01: y = 16'h200;
			16'h3e02: y = 16'h200;
			16'h3e03: y = 16'h200;
			16'h3e04: y = 16'h200;
			16'h3e05: y = 16'h200;
			16'h3e06: y = 16'h200;
			16'h3e07: y = 16'h200;
			16'h3e08: y = 16'h200;
			16'h3e09: y = 16'h200;
			16'h3e0a: y = 16'h200;
			16'h3e0b: y = 16'h200;
			16'h3e0c: y = 16'h200;
			16'h3e0d: y = 16'h200;
			16'h3e0e: y = 16'h200;
			16'h3e0f: y = 16'h200;
			16'h3e10: y = 16'h200;
			16'h3e11: y = 16'h200;
			16'h3e12: y = 16'h200;
			16'h3e13: y = 16'h200;
			16'h3e14: y = 16'h200;
			16'h3e15: y = 16'h200;
			16'h3e16: y = 16'h200;
			16'h3e17: y = 16'h200;
			16'h3e18: y = 16'h200;
			16'h3e19: y = 16'h200;
			16'h3e1a: y = 16'h200;
			16'h3e1b: y = 16'h200;
			16'h3e1c: y = 16'h200;
			16'h3e1d: y = 16'h200;
			16'h3e1e: y = 16'h200;
			16'h3e1f: y = 16'h200;
			16'h3e20: y = 16'h200;
			16'h3e21: y = 16'h200;
			16'h3e22: y = 16'h200;
			16'h3e23: y = 16'h200;
			16'h3e24: y = 16'h200;
			16'h3e25: y = 16'h200;
			16'h3e26: y = 16'h200;
			16'h3e27: y = 16'h200;
			16'h3e28: y = 16'h200;
			16'h3e29: y = 16'h200;
			16'h3e2a: y = 16'h200;
			16'h3e2b: y = 16'h200;
			16'h3e2c: y = 16'h200;
			16'h3e2d: y = 16'h200;
			16'h3e2e: y = 16'h200;
			16'h3e2f: y = 16'h200;
			16'h3e30: y = 16'h200;
			16'h3e31: y = 16'h200;
			16'h3e32: y = 16'h200;
			16'h3e33: y = 16'h200;
			16'h3e34: y = 16'h200;
			16'h3e35: y = 16'h200;
			16'h3e36: y = 16'h200;
			16'h3e37: y = 16'h200;
			16'h3e38: y = 16'h200;
			16'h3e39: y = 16'h200;
			16'h3e3a: y = 16'h200;
			16'h3e3b: y = 16'h200;
			16'h3e3c: y = 16'h200;
			16'h3e3d: y = 16'h200;
			16'h3e3e: y = 16'h200;
			16'h3e3f: y = 16'h200;
			16'h3e40: y = 16'h200;
			16'h3e41: y = 16'h200;
			16'h3e42: y = 16'h200;
			16'h3e43: y = 16'h200;
			16'h3e44: y = 16'h200;
			16'h3e45: y = 16'h200;
			16'h3e46: y = 16'h200;
			16'h3e47: y = 16'h200;
			16'h3e48: y = 16'h200;
			16'h3e49: y = 16'h200;
			16'h3e4a: y = 16'h200;
			16'h3e4b: y = 16'h200;
			16'h3e4c: y = 16'h200;
			16'h3e4d: y = 16'h200;
			16'h3e4e: y = 16'h200;
			16'h3e4f: y = 16'h200;
			16'h3e50: y = 16'h200;
			16'h3e51: y = 16'h200;
			16'h3e52: y = 16'h200;
			16'h3e53: y = 16'h200;
			16'h3e54: y = 16'h200;
			16'h3e55: y = 16'h200;
			16'h3e56: y = 16'h200;
			16'h3e57: y = 16'h200;
			16'h3e58: y = 16'h200;
			16'h3e59: y = 16'h200;
			16'h3e5a: y = 16'h200;
			16'h3e5b: y = 16'h200;
			16'h3e5c: y = 16'h200;
			16'h3e5d: y = 16'h200;
			16'h3e5e: y = 16'h200;
			16'h3e5f: y = 16'h200;
			16'h3e60: y = 16'h200;
			16'h3e61: y = 16'h200;
			16'h3e62: y = 16'h200;
			16'h3e63: y = 16'h200;
			16'h3e64: y = 16'h200;
			16'h3e65: y = 16'h200;
			16'h3e66: y = 16'h200;
			16'h3e67: y = 16'h200;
			16'h3e68: y = 16'h200;
			16'h3e69: y = 16'h200;
			16'h3e6a: y = 16'h200;
			16'h3e6b: y = 16'h200;
			16'h3e6c: y = 16'h200;
			16'h3e6d: y = 16'h200;
			16'h3e6e: y = 16'h200;
			16'h3e6f: y = 16'h200;
			16'h3e70: y = 16'h200;
			16'h3e71: y = 16'h200;
			16'h3e72: y = 16'h200;
			16'h3e73: y = 16'h200;
			16'h3e74: y = 16'h200;
			16'h3e75: y = 16'h200;
			16'h3e76: y = 16'h200;
			16'h3e77: y = 16'h200;
			16'h3e78: y = 16'h200;
			16'h3e79: y = 16'h200;
			16'h3e7a: y = 16'h200;
			16'h3e7b: y = 16'h200;
			16'h3e7c: y = 16'h200;
			16'h3e7d: y = 16'h200;
			16'h3e7e: y = 16'h200;
			16'h3e7f: y = 16'h200;
			16'h3e80: y = 16'h200;
			16'h3e81: y = 16'h200;
			16'h3e82: y = 16'h200;
			16'h3e83: y = 16'h200;
			16'h3e84: y = 16'h200;
			16'h3e85: y = 16'h200;
			16'h3e86: y = 16'h200;
			16'h3e87: y = 16'h200;
			16'h3e88: y = 16'h200;
			16'h3e89: y = 16'h200;
			16'h3e8a: y = 16'h200;
			16'h3e8b: y = 16'h200;
			16'h3e8c: y = 16'h200;
			16'h3e8d: y = 16'h200;
			16'h3e8e: y = 16'h200;
			16'h3e8f: y = 16'h200;
			16'h3e90: y = 16'h200;
			16'h3e91: y = 16'h200;
			16'h3e92: y = 16'h200;
			16'h3e93: y = 16'h200;
			16'h3e94: y = 16'h200;
			16'h3e95: y = 16'h200;
			16'h3e96: y = 16'h200;
			16'h3e97: y = 16'h200;
			16'h3e98: y = 16'h200;
			16'h3e99: y = 16'h200;
			16'h3e9a: y = 16'h200;
			16'h3e9b: y = 16'h200;
			16'h3e9c: y = 16'h200;
			16'h3e9d: y = 16'h200;
			16'h3e9e: y = 16'h200;
			16'h3e9f: y = 16'h200;
			16'h3ea0: y = 16'h200;
			16'h3ea1: y = 16'h200;
			16'h3ea2: y = 16'h200;
			16'h3ea3: y = 16'h200;
			16'h3ea4: y = 16'h200;
			16'h3ea5: y = 16'h200;
			16'h3ea6: y = 16'h200;
			16'h3ea7: y = 16'h200;
			16'h3ea8: y = 16'h200;
			16'h3ea9: y = 16'h200;
			16'h3eaa: y = 16'h200;
			16'h3eab: y = 16'h200;
			16'h3eac: y = 16'h200;
			16'h3ead: y = 16'h200;
			16'h3eae: y = 16'h200;
			16'h3eaf: y = 16'h200;
			16'h3eb0: y = 16'h200;
			16'h3eb1: y = 16'h200;
			16'h3eb2: y = 16'h200;
			16'h3eb3: y = 16'h200;
			16'h3eb4: y = 16'h200;
			16'h3eb5: y = 16'h200;
			16'h3eb6: y = 16'h200;
			16'h3eb7: y = 16'h200;
			16'h3eb8: y = 16'h200;
			16'h3eb9: y = 16'h200;
			16'h3eba: y = 16'h200;
			16'h3ebb: y = 16'h200;
			16'h3ebc: y = 16'h200;
			16'h3ebd: y = 16'h200;
			16'h3ebe: y = 16'h200;
			16'h3ebf: y = 16'h200;
			16'h3ec0: y = 16'h200;
			16'h3ec1: y = 16'h200;
			16'h3ec2: y = 16'h200;
			16'h3ec3: y = 16'h200;
			16'h3ec4: y = 16'h200;
			16'h3ec5: y = 16'h200;
			16'h3ec6: y = 16'h200;
			16'h3ec7: y = 16'h200;
			16'h3ec8: y = 16'h200;
			16'h3ec9: y = 16'h200;
			16'h3eca: y = 16'h200;
			16'h3ecb: y = 16'h200;
			16'h3ecc: y = 16'h200;
			16'h3ecd: y = 16'h200;
			16'h3ece: y = 16'h200;
			16'h3ecf: y = 16'h200;
			16'h3ed0: y = 16'h200;
			16'h3ed1: y = 16'h200;
			16'h3ed2: y = 16'h200;
			16'h3ed3: y = 16'h200;
			16'h3ed4: y = 16'h200;
			16'h3ed5: y = 16'h200;
			16'h3ed6: y = 16'h200;
			16'h3ed7: y = 16'h200;
			16'h3ed8: y = 16'h200;
			16'h3ed9: y = 16'h200;
			16'h3eda: y = 16'h200;
			16'h3edb: y = 16'h200;
			16'h3edc: y = 16'h200;
			16'h3edd: y = 16'h200;
			16'h3ede: y = 16'h200;
			16'h3edf: y = 16'h200;
			16'h3ee0: y = 16'h200;
			16'h3ee1: y = 16'h200;
			16'h3ee2: y = 16'h200;
			16'h3ee3: y = 16'h200;
			16'h3ee4: y = 16'h200;
			16'h3ee5: y = 16'h200;
			16'h3ee6: y = 16'h200;
			16'h3ee7: y = 16'h200;
			16'h3ee8: y = 16'h200;
			16'h3ee9: y = 16'h200;
			16'h3eea: y = 16'h200;
			16'h3eeb: y = 16'h200;
			16'h3eec: y = 16'h200;
			16'h3eed: y = 16'h200;
			16'h3eee: y = 16'h200;
			16'h3eef: y = 16'h200;
			16'h3ef0: y = 16'h200;
			16'h3ef1: y = 16'h200;
			16'h3ef2: y = 16'h200;
			16'h3ef3: y = 16'h200;
			16'h3ef4: y = 16'h200;
			16'h3ef5: y = 16'h200;
			16'h3ef6: y = 16'h200;
			16'h3ef7: y = 16'h200;
			16'h3ef8: y = 16'h200;
			16'h3ef9: y = 16'h200;
			16'h3efa: y = 16'h200;
			16'h3efb: y = 16'h200;
			16'h3efc: y = 16'h200;
			16'h3efd: y = 16'h200;
			16'h3efe: y = 16'h200;
			16'h3eff: y = 16'h200;
			16'h3f00: y = 16'h200;
			16'h3f01: y = 16'h200;
			16'h3f02: y = 16'h200;
			16'h3f03: y = 16'h200;
			16'h3f04: y = 16'h200;
			16'h3f05: y = 16'h200;
			16'h3f06: y = 16'h200;
			16'h3f07: y = 16'h200;
			16'h3f08: y = 16'h200;
			16'h3f09: y = 16'h200;
			16'h3f0a: y = 16'h200;
			16'h3f0b: y = 16'h200;
			16'h3f0c: y = 16'h200;
			16'h3f0d: y = 16'h200;
			16'h3f0e: y = 16'h200;
			16'h3f0f: y = 16'h200;
			16'h3f10: y = 16'h200;
			16'h3f11: y = 16'h200;
			16'h3f12: y = 16'h200;
			16'h3f13: y = 16'h200;
			16'h3f14: y = 16'h200;
			16'h3f15: y = 16'h200;
			16'h3f16: y = 16'h200;
			16'h3f17: y = 16'h200;
			16'h3f18: y = 16'h200;
			16'h3f19: y = 16'h200;
			16'h3f1a: y = 16'h200;
			16'h3f1b: y = 16'h200;
			16'h3f1c: y = 16'h200;
			16'h3f1d: y = 16'h200;
			16'h3f1e: y = 16'h200;
			16'h3f1f: y = 16'h200;
			16'h3f20: y = 16'h200;
			16'h3f21: y = 16'h200;
			16'h3f22: y = 16'h200;
			16'h3f23: y = 16'h200;
			16'h3f24: y = 16'h200;
			16'h3f25: y = 16'h200;
			16'h3f26: y = 16'h200;
			16'h3f27: y = 16'h200;
			16'h3f28: y = 16'h200;
			16'h3f29: y = 16'h200;
			16'h3f2a: y = 16'h200;
			16'h3f2b: y = 16'h200;
			16'h3f2c: y = 16'h200;
			16'h3f2d: y = 16'h200;
			16'h3f2e: y = 16'h200;
			16'h3f2f: y = 16'h200;
			16'h3f30: y = 16'h200;
			16'h3f31: y = 16'h200;
			16'h3f32: y = 16'h200;
			16'h3f33: y = 16'h200;
			16'h3f34: y = 16'h200;
			16'h3f35: y = 16'h200;
			16'h3f36: y = 16'h200;
			16'h3f37: y = 16'h200;
			16'h3f38: y = 16'h200;
			16'h3f39: y = 16'h200;
			16'h3f3a: y = 16'h200;
			16'h3f3b: y = 16'h200;
			16'h3f3c: y = 16'h200;
			16'h3f3d: y = 16'h200;
			16'h3f3e: y = 16'h200;
			16'h3f3f: y = 16'h200;
			16'h3f40: y = 16'h200;
			16'h3f41: y = 16'h200;
			16'h3f42: y = 16'h200;
			16'h3f43: y = 16'h200;
			16'h3f44: y = 16'h200;
			16'h3f45: y = 16'h200;
			16'h3f46: y = 16'h200;
			16'h3f47: y = 16'h200;
			16'h3f48: y = 16'h200;
			16'h3f49: y = 16'h200;
			16'h3f4a: y = 16'h200;
			16'h3f4b: y = 16'h200;
			16'h3f4c: y = 16'h200;
			16'h3f4d: y = 16'h200;
			16'h3f4e: y = 16'h200;
			16'h3f4f: y = 16'h200;
			16'h3f50: y = 16'h200;
			16'h3f51: y = 16'h200;
			16'h3f52: y = 16'h200;
			16'h3f53: y = 16'h200;
			16'h3f54: y = 16'h200;
			16'h3f55: y = 16'h200;
			16'h3f56: y = 16'h200;
			16'h3f57: y = 16'h200;
			16'h3f58: y = 16'h200;
			16'h3f59: y = 16'h200;
			16'h3f5a: y = 16'h200;
			16'h3f5b: y = 16'h200;
			16'h3f5c: y = 16'h200;
			16'h3f5d: y = 16'h200;
			16'h3f5e: y = 16'h200;
			16'h3f5f: y = 16'h200;
			16'h3f60: y = 16'h200;
			16'h3f61: y = 16'h200;
			16'h3f62: y = 16'h200;
			16'h3f63: y = 16'h200;
			16'h3f64: y = 16'h200;
			16'h3f65: y = 16'h200;
			16'h3f66: y = 16'h200;
			16'h3f67: y = 16'h200;
			16'h3f68: y = 16'h200;
			16'h3f69: y = 16'h200;
			16'h3f6a: y = 16'h200;
			16'h3f6b: y = 16'h200;
			16'h3f6c: y = 16'h200;
			16'h3f6d: y = 16'h200;
			16'h3f6e: y = 16'h200;
			16'h3f6f: y = 16'h200;
			16'h3f70: y = 16'h200;
			16'h3f71: y = 16'h200;
			16'h3f72: y = 16'h200;
			16'h3f73: y = 16'h200;
			16'h3f74: y = 16'h200;
			16'h3f75: y = 16'h200;
			16'h3f76: y = 16'h200;
			16'h3f77: y = 16'h200;
			16'h3f78: y = 16'h200;
			16'h3f79: y = 16'h200;
			16'h3f7a: y = 16'h200;
			16'h3f7b: y = 16'h200;
			16'h3f7c: y = 16'h200;
			16'h3f7d: y = 16'h200;
			16'h3f7e: y = 16'h200;
			16'h3f7f: y = 16'h200;
			16'h3f80: y = 16'h200;
			16'h3f81: y = 16'h200;
			16'h3f82: y = 16'h200;
			16'h3f83: y = 16'h200;
			16'h3f84: y = 16'h200;
			16'h3f85: y = 16'h200;
			16'h3f86: y = 16'h200;
			16'h3f87: y = 16'h200;
			16'h3f88: y = 16'h200;
			16'h3f89: y = 16'h200;
			16'h3f8a: y = 16'h200;
			16'h3f8b: y = 16'h200;
			16'h3f8c: y = 16'h200;
			16'h3f8d: y = 16'h200;
			16'h3f8e: y = 16'h200;
			16'h3f8f: y = 16'h200;
			16'h3f90: y = 16'h200;
			16'h3f91: y = 16'h200;
			16'h3f92: y = 16'h200;
			16'h3f93: y = 16'h200;
			16'h3f94: y = 16'h200;
			16'h3f95: y = 16'h200;
			16'h3f96: y = 16'h200;
			16'h3f97: y = 16'h200;
			16'h3f98: y = 16'h200;
			16'h3f99: y = 16'h200;
			16'h3f9a: y = 16'h200;
			16'h3f9b: y = 16'h200;
			16'h3f9c: y = 16'h200;
			16'h3f9d: y = 16'h200;
			16'h3f9e: y = 16'h200;
			16'h3f9f: y = 16'h200;
			16'h3fa0: y = 16'h200;
			16'h3fa1: y = 16'h200;
			16'h3fa2: y = 16'h200;
			16'h3fa3: y = 16'h200;
			16'h3fa4: y = 16'h200;
			16'h3fa5: y = 16'h200;
			16'h3fa6: y = 16'h200;
			16'h3fa7: y = 16'h200;
			16'h3fa8: y = 16'h200;
			16'h3fa9: y = 16'h200;
			16'h3faa: y = 16'h200;
			16'h3fab: y = 16'h200;
			16'h3fac: y = 16'h200;
			16'h3fad: y = 16'h200;
			16'h3fae: y = 16'h200;
			16'h3faf: y = 16'h200;
			16'h3fb0: y = 16'h200;
			16'h3fb1: y = 16'h200;
			16'h3fb2: y = 16'h200;
			16'h3fb3: y = 16'h200;
			16'h3fb4: y = 16'h200;
			16'h3fb5: y = 16'h200;
			16'h3fb6: y = 16'h200;
			16'h3fb7: y = 16'h200;
			16'h3fb8: y = 16'h200;
			16'h3fb9: y = 16'h200;
			16'h3fba: y = 16'h200;
			16'h3fbb: y = 16'h200;
			16'h3fbc: y = 16'h200;
			16'h3fbd: y = 16'h200;
			16'h3fbe: y = 16'h200;
			16'h3fbf: y = 16'h200;
			16'h3fc0: y = 16'h200;
			16'h3fc1: y = 16'h200;
			16'h3fc2: y = 16'h200;
			16'h3fc3: y = 16'h200;
			16'h3fc4: y = 16'h200;
			16'h3fc5: y = 16'h200;
			16'h3fc6: y = 16'h200;
			16'h3fc7: y = 16'h200;
			16'h3fc8: y = 16'h200;
			16'h3fc9: y = 16'h200;
			16'h3fca: y = 16'h200;
			16'h3fcb: y = 16'h200;
			16'h3fcc: y = 16'h200;
			16'h3fcd: y = 16'h200;
			16'h3fce: y = 16'h200;
			16'h3fcf: y = 16'h200;
			16'h3fd0: y = 16'h200;
			16'h3fd1: y = 16'h200;
			16'h3fd2: y = 16'h200;
			16'h3fd3: y = 16'h200;
			16'h3fd4: y = 16'h200;
			16'h3fd5: y = 16'h200;
			16'h3fd6: y = 16'h200;
			16'h3fd7: y = 16'h200;
			16'h3fd8: y = 16'h200;
			16'h3fd9: y = 16'h200;
			16'h3fda: y = 16'h200;
			16'h3fdb: y = 16'h200;
			16'h3fdc: y = 16'h200;
			16'h3fdd: y = 16'h200;
			16'h3fde: y = 16'h200;
			16'h3fdf: y = 16'h200;
			16'h3fe0: y = 16'h200;
			16'h3fe1: y = 16'h200;
			16'h3fe2: y = 16'h200;
			16'h3fe3: y = 16'h200;
			16'h3fe4: y = 16'h200;
			16'h3fe5: y = 16'h200;
			16'h3fe6: y = 16'h200;
			16'h3fe7: y = 16'h200;
			16'h3fe8: y = 16'h200;
			16'h3fe9: y = 16'h200;
			16'h3fea: y = 16'h200;
			16'h3feb: y = 16'h200;
			16'h3fec: y = 16'h200;
			16'h3fed: y = 16'h200;
			16'h3fee: y = 16'h200;
			16'h3fef: y = 16'h200;
			16'h3ff0: y = 16'h200;
			16'h3ff1: y = 16'h200;
			16'h3ff2: y = 16'h200;
			16'h3ff3: y = 16'h200;
			16'h3ff4: y = 16'h200;
			16'h3ff5: y = 16'h200;
			16'h3ff6: y = 16'h200;
			16'h3ff7: y = 16'h200;
			16'h3ff8: y = 16'h200;
			16'h3ff9: y = 16'h200;
			16'h3ffa: y = 16'h200;
			16'h3ffb: y = 16'h200;
			16'h3ffc: y = 16'h200;
			16'h3ffd: y = 16'h200;
			16'h3ffe: y = 16'h200;
			16'h3fff: y = 16'h200;
			16'h4000: y = 16'h200;
			16'h4001: y = 16'h200;
			16'h4002: y = 16'h200;
			16'h4003: y = 16'h200;
			16'h4004: y = 16'h200;
			16'h4005: y = 16'h200;
			16'h4006: y = 16'h200;
			16'h4007: y = 16'h200;
			16'h4008: y = 16'h200;
			16'h4009: y = 16'h200;
			16'h400a: y = 16'h200;
			16'h400b: y = 16'h200;
			16'h400c: y = 16'h200;
			16'h400d: y = 16'h200;
			16'h400e: y = 16'h200;
			16'h400f: y = 16'h200;
			16'h4010: y = 16'h200;
			16'h4011: y = 16'h200;
			16'h4012: y = 16'h200;
			16'h4013: y = 16'h200;
			16'h4014: y = 16'h200;
			16'h4015: y = 16'h200;
			16'h4016: y = 16'h200;
			16'h4017: y = 16'h200;
			16'h4018: y = 16'h200;
			16'h4019: y = 16'h200;
			16'h401a: y = 16'h200;
			16'h401b: y = 16'h200;
			16'h401c: y = 16'h200;
			16'h401d: y = 16'h200;
			16'h401e: y = 16'h200;
			16'h401f: y = 16'h200;
			16'h4020: y = 16'h200;
			16'h4021: y = 16'h200;
			16'h4022: y = 16'h200;
			16'h4023: y = 16'h200;
			16'h4024: y = 16'h200;
			16'h4025: y = 16'h200;
			16'h4026: y = 16'h200;
			16'h4027: y = 16'h200;
			16'h4028: y = 16'h200;
			16'h4029: y = 16'h200;
			16'h402a: y = 16'h200;
			16'h402b: y = 16'h200;
			16'h402c: y = 16'h200;
			16'h402d: y = 16'h200;
			16'h402e: y = 16'h200;
			16'h402f: y = 16'h200;
			16'h4030: y = 16'h200;
			16'h4031: y = 16'h200;
			16'h4032: y = 16'h200;
			16'h4033: y = 16'h200;
			16'h4034: y = 16'h200;
			16'h4035: y = 16'h200;
			16'h4036: y = 16'h200;
			16'h4037: y = 16'h200;
			16'h4038: y = 16'h200;
			16'h4039: y = 16'h200;
			16'h403a: y = 16'h200;
			16'h403b: y = 16'h200;
			16'h403c: y = 16'h200;
			16'h403d: y = 16'h200;
			16'h403e: y = 16'h200;
			16'h403f: y = 16'h200;
			16'h4040: y = 16'h200;
			16'h4041: y = 16'h200;
			16'h4042: y = 16'h200;
			16'h4043: y = 16'h200;
			16'h4044: y = 16'h200;
			16'h4045: y = 16'h200;
			16'h4046: y = 16'h200;
			16'h4047: y = 16'h200;
			16'h4048: y = 16'h200;
			16'h4049: y = 16'h200;
			16'h404a: y = 16'h200;
			16'h404b: y = 16'h200;
			16'h404c: y = 16'h200;
			16'h404d: y = 16'h200;
			16'h404e: y = 16'h200;
			16'h404f: y = 16'h200;
			16'h4050: y = 16'h200;
			16'h4051: y = 16'h200;
			16'h4052: y = 16'h200;
			16'h4053: y = 16'h200;
			16'h4054: y = 16'h200;
			16'h4055: y = 16'h200;
			16'h4056: y = 16'h200;
			16'h4057: y = 16'h200;
			16'h4058: y = 16'h200;
			16'h4059: y = 16'h200;
			16'h405a: y = 16'h200;
			16'h405b: y = 16'h200;
			16'h405c: y = 16'h200;
			16'h405d: y = 16'h200;
			16'h405e: y = 16'h200;
			16'h405f: y = 16'h200;
			16'h4060: y = 16'h200;
			16'h4061: y = 16'h200;
			16'h4062: y = 16'h200;
			16'h4063: y = 16'h200;
			16'h4064: y = 16'h200;
			16'h4065: y = 16'h200;
			16'h4066: y = 16'h200;
			16'h4067: y = 16'h200;
			16'h4068: y = 16'h200;
			16'h4069: y = 16'h200;
			16'h406a: y = 16'h200;
			16'h406b: y = 16'h200;
			16'h406c: y = 16'h200;
			16'h406d: y = 16'h200;
			16'h406e: y = 16'h200;
			16'h406f: y = 16'h200;
			16'h4070: y = 16'h200;
			16'h4071: y = 16'h200;
			16'h4072: y = 16'h200;
			16'h4073: y = 16'h200;
			16'h4074: y = 16'h200;
			16'h4075: y = 16'h200;
			16'h4076: y = 16'h200;
			16'h4077: y = 16'h200;
			16'h4078: y = 16'h200;
			16'h4079: y = 16'h200;
			16'h407a: y = 16'h200;
			16'h407b: y = 16'h200;
			16'h407c: y = 16'h200;
			16'h407d: y = 16'h200;
			16'h407e: y = 16'h200;
			16'h407f: y = 16'h200;
			16'h4080: y = 16'h200;
			16'h4081: y = 16'h200;
			16'h4082: y = 16'h200;
			16'h4083: y = 16'h200;
			16'h4084: y = 16'h200;
			16'h4085: y = 16'h200;
			16'h4086: y = 16'h200;
			16'h4087: y = 16'h200;
			16'h4088: y = 16'h200;
			16'h4089: y = 16'h200;
			16'h408a: y = 16'h200;
			16'h408b: y = 16'h200;
			16'h408c: y = 16'h200;
			16'h408d: y = 16'h200;
			16'h408e: y = 16'h200;
			16'h408f: y = 16'h200;
			16'h4090: y = 16'h200;
			16'h4091: y = 16'h200;
			16'h4092: y = 16'h200;
			16'h4093: y = 16'h200;
			16'h4094: y = 16'h200;
			16'h4095: y = 16'h200;
			16'h4096: y = 16'h200;
			16'h4097: y = 16'h200;
			16'h4098: y = 16'h200;
			16'h4099: y = 16'h200;
			16'h409a: y = 16'h200;
			16'h409b: y = 16'h200;
			16'h409c: y = 16'h200;
			16'h409d: y = 16'h200;
			16'h409e: y = 16'h200;
			16'h409f: y = 16'h200;
			16'h40a0: y = 16'h200;
			16'h40a1: y = 16'h200;
			16'h40a2: y = 16'h200;
			16'h40a3: y = 16'h200;
			16'h40a4: y = 16'h200;
			16'h40a5: y = 16'h200;
			16'h40a6: y = 16'h200;
			16'h40a7: y = 16'h200;
			16'h40a8: y = 16'h200;
			16'h40a9: y = 16'h200;
			16'h40aa: y = 16'h200;
			16'h40ab: y = 16'h200;
			16'h40ac: y = 16'h200;
			16'h40ad: y = 16'h200;
			16'h40ae: y = 16'h200;
			16'h40af: y = 16'h200;
			16'h40b0: y = 16'h200;
			16'h40b1: y = 16'h200;
			16'h40b2: y = 16'h200;
			16'h40b3: y = 16'h200;
			16'h40b4: y = 16'h200;
			16'h40b5: y = 16'h200;
			16'h40b6: y = 16'h200;
			16'h40b7: y = 16'h200;
			16'h40b8: y = 16'h200;
			16'h40b9: y = 16'h200;
			16'h40ba: y = 16'h200;
			16'h40bb: y = 16'h200;
			16'h40bc: y = 16'h200;
			16'h40bd: y = 16'h200;
			16'h40be: y = 16'h200;
			16'h40bf: y = 16'h200;
			16'h40c0: y = 16'h200;
			16'h40c1: y = 16'h200;
			16'h40c2: y = 16'h200;
			16'h40c3: y = 16'h200;
			16'h40c4: y = 16'h200;
			16'h40c5: y = 16'h200;
			16'h40c6: y = 16'h200;
			16'h40c7: y = 16'h200;
			16'h40c8: y = 16'h200;
			16'h40c9: y = 16'h200;
			16'h40ca: y = 16'h200;
			16'h40cb: y = 16'h200;
			16'h40cc: y = 16'h200;
			16'h40cd: y = 16'h200;
			16'h40ce: y = 16'h200;
			16'h40cf: y = 16'h200;
			16'h40d0: y = 16'h200;
			16'h40d1: y = 16'h200;
			16'h40d2: y = 16'h200;
			16'h40d3: y = 16'h200;
			16'h40d4: y = 16'h200;
			16'h40d5: y = 16'h200;
			16'h40d6: y = 16'h200;
			16'h40d7: y = 16'h200;
			16'h40d8: y = 16'h200;
			16'h40d9: y = 16'h200;
			16'h40da: y = 16'h200;
			16'h40db: y = 16'h200;
			16'h40dc: y = 16'h200;
			16'h40dd: y = 16'h200;
			16'h40de: y = 16'h200;
			16'h40df: y = 16'h200;
			16'h40e0: y = 16'h200;
			16'h40e1: y = 16'h200;
			16'h40e2: y = 16'h200;
			16'h40e3: y = 16'h200;
			16'h40e4: y = 16'h200;
			16'h40e5: y = 16'h200;
			16'h40e6: y = 16'h200;
			16'h40e7: y = 16'h200;
			16'h40e8: y = 16'h200;
			16'h40e9: y = 16'h200;
			16'h40ea: y = 16'h200;
			16'h40eb: y = 16'h200;
			16'h40ec: y = 16'h200;
			16'h40ed: y = 16'h200;
			16'h40ee: y = 16'h200;
			16'h40ef: y = 16'h200;
			16'h40f0: y = 16'h200;
			16'h40f1: y = 16'h200;
			16'h40f2: y = 16'h200;
			16'h40f3: y = 16'h200;
			16'h40f4: y = 16'h200;
			16'h40f5: y = 16'h200;
			16'h40f6: y = 16'h200;
			16'h40f7: y = 16'h200;
			16'h40f8: y = 16'h200;
			16'h40f9: y = 16'h200;
			16'h40fa: y = 16'h200;
			16'h40fb: y = 16'h200;
			16'h40fc: y = 16'h200;
			16'h40fd: y = 16'h200;
			16'h40fe: y = 16'h200;
			16'h40ff: y = 16'h200;
			16'h4100: y = 16'h200;
			16'h4101: y = 16'h200;
			16'h4102: y = 16'h200;
			16'h4103: y = 16'h200;
			16'h4104: y = 16'h200;
			16'h4105: y = 16'h200;
			16'h4106: y = 16'h200;
			16'h4107: y = 16'h200;
			16'h4108: y = 16'h200;
			16'h4109: y = 16'h200;
			16'h410a: y = 16'h200;
			16'h410b: y = 16'h200;
			16'h410c: y = 16'h200;
			16'h410d: y = 16'h200;
			16'h410e: y = 16'h200;
			16'h410f: y = 16'h200;
			16'h4110: y = 16'h200;
			16'h4111: y = 16'h200;
			16'h4112: y = 16'h200;
			16'h4113: y = 16'h200;
			16'h4114: y = 16'h200;
			16'h4115: y = 16'h200;
			16'h4116: y = 16'h200;
			16'h4117: y = 16'h200;
			16'h4118: y = 16'h200;
			16'h4119: y = 16'h200;
			16'h411a: y = 16'h200;
			16'h411b: y = 16'h200;
			16'h411c: y = 16'h200;
			16'h411d: y = 16'h200;
			16'h411e: y = 16'h200;
			16'h411f: y = 16'h200;
			16'h4120: y = 16'h200;
			16'h4121: y = 16'h200;
			16'h4122: y = 16'h200;
			16'h4123: y = 16'h200;
			16'h4124: y = 16'h200;
			16'h4125: y = 16'h200;
			16'h4126: y = 16'h200;
			16'h4127: y = 16'h200;
			16'h4128: y = 16'h200;
			16'h4129: y = 16'h200;
			16'h412a: y = 16'h200;
			16'h412b: y = 16'h200;
			16'h412c: y = 16'h200;
			16'h412d: y = 16'h200;
			16'h412e: y = 16'h200;
			16'h412f: y = 16'h200;
			16'h4130: y = 16'h200;
			16'h4131: y = 16'h200;
			16'h4132: y = 16'h200;
			16'h4133: y = 16'h200;
			16'h4134: y = 16'h200;
			16'h4135: y = 16'h200;
			16'h4136: y = 16'h200;
			16'h4137: y = 16'h200;
			16'h4138: y = 16'h200;
			16'h4139: y = 16'h200;
			16'h413a: y = 16'h200;
			16'h413b: y = 16'h200;
			16'h413c: y = 16'h200;
			16'h413d: y = 16'h200;
			16'h413e: y = 16'h200;
			16'h413f: y = 16'h200;
			16'h4140: y = 16'h200;
			16'h4141: y = 16'h200;
			16'h4142: y = 16'h200;
			16'h4143: y = 16'h200;
			16'h4144: y = 16'h200;
			16'h4145: y = 16'h200;
			16'h4146: y = 16'h200;
			16'h4147: y = 16'h200;
			16'h4148: y = 16'h200;
			16'h4149: y = 16'h200;
			16'h414a: y = 16'h200;
			16'h414b: y = 16'h200;
			16'h414c: y = 16'h200;
			16'h414d: y = 16'h200;
			16'h414e: y = 16'h200;
			16'h414f: y = 16'h200;
			16'h4150: y = 16'h200;
			16'h4151: y = 16'h200;
			16'h4152: y = 16'h200;
			16'h4153: y = 16'h200;
			16'h4154: y = 16'h200;
			16'h4155: y = 16'h200;
			16'h4156: y = 16'h200;
			16'h4157: y = 16'h200;
			16'h4158: y = 16'h200;
			16'h4159: y = 16'h200;
			16'h415a: y = 16'h200;
			16'h415b: y = 16'h200;
			16'h415c: y = 16'h200;
			16'h415d: y = 16'h200;
			16'h415e: y = 16'h200;
			16'h415f: y = 16'h200;
			16'h4160: y = 16'h200;
			16'h4161: y = 16'h200;
			16'h4162: y = 16'h200;
			16'h4163: y = 16'h200;
			16'h4164: y = 16'h200;
			16'h4165: y = 16'h200;
			16'h4166: y = 16'h200;
			16'h4167: y = 16'h200;
			16'h4168: y = 16'h200;
			16'h4169: y = 16'h200;
			16'h416a: y = 16'h200;
			16'h416b: y = 16'h200;
			16'h416c: y = 16'h200;
			16'h416d: y = 16'h200;
			16'h416e: y = 16'h200;
			16'h416f: y = 16'h200;
			16'h4170: y = 16'h200;
			16'h4171: y = 16'h200;
			16'h4172: y = 16'h200;
			16'h4173: y = 16'h200;
			16'h4174: y = 16'h200;
			16'h4175: y = 16'h200;
			16'h4176: y = 16'h200;
			16'h4177: y = 16'h200;
			16'h4178: y = 16'h200;
			16'h4179: y = 16'h200;
			16'h417a: y = 16'h200;
			16'h417b: y = 16'h200;
			16'h417c: y = 16'h200;
			16'h417d: y = 16'h200;
			16'h417e: y = 16'h200;
			16'h417f: y = 16'h200;
			16'h4180: y = 16'h200;
			16'h4181: y = 16'h200;
			16'h4182: y = 16'h200;
			16'h4183: y = 16'h200;
			16'h4184: y = 16'h200;
			16'h4185: y = 16'h200;
			16'h4186: y = 16'h200;
			16'h4187: y = 16'h200;
			16'h4188: y = 16'h200;
			16'h4189: y = 16'h200;
			16'h418a: y = 16'h200;
			16'h418b: y = 16'h200;
			16'h418c: y = 16'h200;
			16'h418d: y = 16'h200;
			16'h418e: y = 16'h200;
			16'h418f: y = 16'h200;
			16'h4190: y = 16'h200;
			16'h4191: y = 16'h200;
			16'h4192: y = 16'h200;
			16'h4193: y = 16'h200;
			16'h4194: y = 16'h200;
			16'h4195: y = 16'h200;
			16'h4196: y = 16'h200;
			16'h4197: y = 16'h200;
			16'h4198: y = 16'h200;
			16'h4199: y = 16'h200;
			16'h419a: y = 16'h200;
			16'h419b: y = 16'h200;
			16'h419c: y = 16'h200;
			16'h419d: y = 16'h200;
			16'h419e: y = 16'h200;
			16'h419f: y = 16'h200;
			16'h41a0: y = 16'h200;
			16'h41a1: y = 16'h200;
			16'h41a2: y = 16'h200;
			16'h41a3: y = 16'h200;
			16'h41a4: y = 16'h200;
			16'h41a5: y = 16'h200;
			16'h41a6: y = 16'h200;
			16'h41a7: y = 16'h200;
			16'h41a8: y = 16'h200;
			16'h41a9: y = 16'h200;
			16'h41aa: y = 16'h200;
			16'h41ab: y = 16'h200;
			16'h41ac: y = 16'h200;
			16'h41ad: y = 16'h200;
			16'h41ae: y = 16'h200;
			16'h41af: y = 16'h200;
			16'h41b0: y = 16'h200;
			16'h41b1: y = 16'h200;
			16'h41b2: y = 16'h200;
			16'h41b3: y = 16'h200;
			16'h41b4: y = 16'h200;
			16'h41b5: y = 16'h200;
			16'h41b6: y = 16'h200;
			16'h41b7: y = 16'h200;
			16'h41b8: y = 16'h200;
			16'h41b9: y = 16'h200;
			16'h41ba: y = 16'h200;
			16'h41bb: y = 16'h200;
			16'h41bc: y = 16'h200;
			16'h41bd: y = 16'h200;
			16'h41be: y = 16'h200;
			16'h41bf: y = 16'h200;
			16'h41c0: y = 16'h200;
			16'h41c1: y = 16'h200;
			16'h41c2: y = 16'h200;
			16'h41c3: y = 16'h200;
			16'h41c4: y = 16'h200;
			16'h41c5: y = 16'h200;
			16'h41c6: y = 16'h200;
			16'h41c7: y = 16'h200;
			16'h41c8: y = 16'h200;
			16'h41c9: y = 16'h200;
			16'h41ca: y = 16'h200;
			16'h41cb: y = 16'h200;
			16'h41cc: y = 16'h200;
			16'h41cd: y = 16'h200;
			16'h41ce: y = 16'h200;
			16'h41cf: y = 16'h200;
			16'h41d0: y = 16'h200;
			16'h41d1: y = 16'h200;
			16'h41d2: y = 16'h200;
			16'h41d3: y = 16'h200;
			16'h41d4: y = 16'h200;
			16'h41d5: y = 16'h200;
			16'h41d6: y = 16'h200;
			16'h41d7: y = 16'h200;
			16'h41d8: y = 16'h200;
			16'h41d9: y = 16'h200;
			16'h41da: y = 16'h200;
			16'h41db: y = 16'h200;
			16'h41dc: y = 16'h200;
			16'h41dd: y = 16'h200;
			16'h41de: y = 16'h200;
			16'h41df: y = 16'h200;
			16'h41e0: y = 16'h200;
			16'h41e1: y = 16'h200;
			16'h41e2: y = 16'h200;
			16'h41e3: y = 16'h200;
			16'h41e4: y = 16'h200;
			16'h41e5: y = 16'h200;
			16'h41e6: y = 16'h200;
			16'h41e7: y = 16'h200;
			16'h41e8: y = 16'h200;
			16'h41e9: y = 16'h200;
			16'h41ea: y = 16'h200;
			16'h41eb: y = 16'h200;
			16'h41ec: y = 16'h200;
			16'h41ed: y = 16'h200;
			16'h41ee: y = 16'h200;
			16'h41ef: y = 16'h200;
			16'h41f0: y = 16'h200;
			16'h41f1: y = 16'h200;
			16'h41f2: y = 16'h200;
			16'h41f3: y = 16'h200;
			16'h41f4: y = 16'h200;
			16'h41f5: y = 16'h200;
			16'h41f6: y = 16'h200;
			16'h41f7: y = 16'h200;
			16'h41f8: y = 16'h200;
			16'h41f9: y = 16'h200;
			16'h41fa: y = 16'h200;
			16'h41fb: y = 16'h200;
			16'h41fc: y = 16'h200;
			16'h41fd: y = 16'h200;
			16'h41fe: y = 16'h200;
			16'h41ff: y = 16'h200;
			16'h4200: y = 16'h200;
			16'h4201: y = 16'h200;
			16'h4202: y = 16'h200;
			16'h4203: y = 16'h200;
			16'h4204: y = 16'h200;
			16'h4205: y = 16'h200;
			16'h4206: y = 16'h200;
			16'h4207: y = 16'h200;
			16'h4208: y = 16'h200;
			16'h4209: y = 16'h200;
			16'h420a: y = 16'h200;
			16'h420b: y = 16'h200;
			16'h420c: y = 16'h200;
			16'h420d: y = 16'h200;
			16'h420e: y = 16'h200;
			16'h420f: y = 16'h200;
			16'h4210: y = 16'h200;
			16'h4211: y = 16'h200;
			16'h4212: y = 16'h200;
			16'h4213: y = 16'h200;
			16'h4214: y = 16'h200;
			16'h4215: y = 16'h200;
			16'h4216: y = 16'h200;
			16'h4217: y = 16'h200;
			16'h4218: y = 16'h200;
			16'h4219: y = 16'h200;
			16'h421a: y = 16'h200;
			16'h421b: y = 16'h200;
			16'h421c: y = 16'h200;
			16'h421d: y = 16'h200;
			16'h421e: y = 16'h200;
			16'h421f: y = 16'h200;
			16'h4220: y = 16'h200;
			16'h4221: y = 16'h200;
			16'h4222: y = 16'h200;
			16'h4223: y = 16'h200;
			16'h4224: y = 16'h200;
			16'h4225: y = 16'h200;
			16'h4226: y = 16'h200;
			16'h4227: y = 16'h200;
			16'h4228: y = 16'h200;
			16'h4229: y = 16'h200;
			16'h422a: y = 16'h200;
			16'h422b: y = 16'h200;
			16'h422c: y = 16'h200;
			16'h422d: y = 16'h200;
			16'h422e: y = 16'h200;
			16'h422f: y = 16'h200;
			16'h4230: y = 16'h200;
			16'h4231: y = 16'h200;
			16'h4232: y = 16'h200;
			16'h4233: y = 16'h200;
			16'h4234: y = 16'h200;
			16'h4235: y = 16'h200;
			16'h4236: y = 16'h200;
			16'h4237: y = 16'h200;
			16'h4238: y = 16'h200;
			16'h4239: y = 16'h200;
			16'h423a: y = 16'h200;
			16'h423b: y = 16'h200;
			16'h423c: y = 16'h200;
			16'h423d: y = 16'h200;
			16'h423e: y = 16'h200;
			16'h423f: y = 16'h200;
			16'h4240: y = 16'h200;
			16'h4241: y = 16'h200;
			16'h4242: y = 16'h200;
			16'h4243: y = 16'h200;
			16'h4244: y = 16'h200;
			16'h4245: y = 16'h200;
			16'h4246: y = 16'h200;
			16'h4247: y = 16'h200;
			16'h4248: y = 16'h200;
			16'h4249: y = 16'h200;
			16'h424a: y = 16'h200;
			16'h424b: y = 16'h200;
			16'h424c: y = 16'h200;
			16'h424d: y = 16'h200;
			16'h424e: y = 16'h200;
			16'h424f: y = 16'h200;
			16'h4250: y = 16'h200;
			16'h4251: y = 16'h200;
			16'h4252: y = 16'h200;
			16'h4253: y = 16'h200;
			16'h4254: y = 16'h200;
			16'h4255: y = 16'h200;
			16'h4256: y = 16'h200;
			16'h4257: y = 16'h200;
			16'h4258: y = 16'h200;
			16'h4259: y = 16'h200;
			16'h425a: y = 16'h200;
			16'h425b: y = 16'h200;
			16'h425c: y = 16'h200;
			16'h425d: y = 16'h200;
			16'h425e: y = 16'h200;
			16'h425f: y = 16'h200;
			16'h4260: y = 16'h200;
			16'h4261: y = 16'h200;
			16'h4262: y = 16'h200;
			16'h4263: y = 16'h200;
			16'h4264: y = 16'h200;
			16'h4265: y = 16'h200;
			16'h4266: y = 16'h200;
			16'h4267: y = 16'h200;
			16'h4268: y = 16'h200;
			16'h4269: y = 16'h200;
			16'h426a: y = 16'h200;
			16'h426b: y = 16'h200;
			16'h426c: y = 16'h200;
			16'h426d: y = 16'h200;
			16'h426e: y = 16'h200;
			16'h426f: y = 16'h200;
			16'h4270: y = 16'h200;
			16'h4271: y = 16'h200;
			16'h4272: y = 16'h200;
			16'h4273: y = 16'h200;
			16'h4274: y = 16'h200;
			16'h4275: y = 16'h200;
			16'h4276: y = 16'h200;
			16'h4277: y = 16'h200;
			16'h4278: y = 16'h200;
			16'h4279: y = 16'h200;
			16'h427a: y = 16'h200;
			16'h427b: y = 16'h200;
			16'h427c: y = 16'h200;
			16'h427d: y = 16'h200;
			16'h427e: y = 16'h200;
			16'h427f: y = 16'h200;
			16'h4280: y = 16'h200;
			16'h4281: y = 16'h200;
			16'h4282: y = 16'h200;
			16'h4283: y = 16'h200;
			16'h4284: y = 16'h200;
			16'h4285: y = 16'h200;
			16'h4286: y = 16'h200;
			16'h4287: y = 16'h200;
			16'h4288: y = 16'h200;
			16'h4289: y = 16'h200;
			16'h428a: y = 16'h200;
			16'h428b: y = 16'h200;
			16'h428c: y = 16'h200;
			16'h428d: y = 16'h200;
			16'h428e: y = 16'h200;
			16'h428f: y = 16'h200;
			16'h4290: y = 16'h200;
			16'h4291: y = 16'h200;
			16'h4292: y = 16'h200;
			16'h4293: y = 16'h200;
			16'h4294: y = 16'h200;
			16'h4295: y = 16'h200;
			16'h4296: y = 16'h200;
			16'h4297: y = 16'h200;
			16'h4298: y = 16'h200;
			16'h4299: y = 16'h200;
			16'h429a: y = 16'h200;
			16'h429b: y = 16'h200;
			16'h429c: y = 16'h200;
			16'h429d: y = 16'h200;
			16'h429e: y = 16'h200;
			16'h429f: y = 16'h200;
			16'h42a0: y = 16'h200;
			16'h42a1: y = 16'h200;
			16'h42a2: y = 16'h200;
			16'h42a3: y = 16'h200;
			16'h42a4: y = 16'h200;
			16'h42a5: y = 16'h200;
			16'h42a6: y = 16'h200;
			16'h42a7: y = 16'h200;
			16'h42a8: y = 16'h200;
			16'h42a9: y = 16'h200;
			16'h42aa: y = 16'h200;
			16'h42ab: y = 16'h200;
			16'h42ac: y = 16'h200;
			16'h42ad: y = 16'h200;
			16'h42ae: y = 16'h200;
			16'h42af: y = 16'h200;
			16'h42b0: y = 16'h200;
			16'h42b1: y = 16'h200;
			16'h42b2: y = 16'h200;
			16'h42b3: y = 16'h200;
			16'h42b4: y = 16'h200;
			16'h42b5: y = 16'h200;
			16'h42b6: y = 16'h200;
			16'h42b7: y = 16'h200;
			16'h42b8: y = 16'h200;
			16'h42b9: y = 16'h200;
			16'h42ba: y = 16'h200;
			16'h42bb: y = 16'h200;
			16'h42bc: y = 16'h200;
			16'h42bd: y = 16'h200;
			16'h42be: y = 16'h200;
			16'h42bf: y = 16'h200;
			16'h42c0: y = 16'h200;
			16'h42c1: y = 16'h200;
			16'h42c2: y = 16'h200;
			16'h42c3: y = 16'h200;
			16'h42c4: y = 16'h200;
			16'h42c5: y = 16'h200;
			16'h42c6: y = 16'h200;
			16'h42c7: y = 16'h200;
			16'h42c8: y = 16'h200;
			16'h42c9: y = 16'h200;
			16'h42ca: y = 16'h200;
			16'h42cb: y = 16'h200;
			16'h42cc: y = 16'h200;
			16'h42cd: y = 16'h200;
			16'h42ce: y = 16'h200;
			16'h42cf: y = 16'h200;
			16'h42d0: y = 16'h200;
			16'h42d1: y = 16'h200;
			16'h42d2: y = 16'h200;
			16'h42d3: y = 16'h200;
			16'h42d4: y = 16'h200;
			16'h42d5: y = 16'h200;
			16'h42d6: y = 16'h200;
			16'h42d7: y = 16'h200;
			16'h42d8: y = 16'h200;
			16'h42d9: y = 16'h200;
			16'h42da: y = 16'h200;
			16'h42db: y = 16'h200;
			16'h42dc: y = 16'h200;
			16'h42dd: y = 16'h200;
			16'h42de: y = 16'h200;
			16'h42df: y = 16'h200;
			16'h42e0: y = 16'h200;
			16'h42e1: y = 16'h200;
			16'h42e2: y = 16'h200;
			16'h42e3: y = 16'h200;
			16'h42e4: y = 16'h200;
			16'h42e5: y = 16'h200;
			16'h42e6: y = 16'h200;
			16'h42e7: y = 16'h200;
			16'h42e8: y = 16'h200;
			16'h42e9: y = 16'h200;
			16'h42ea: y = 16'h200;
			16'h42eb: y = 16'h200;
			16'h42ec: y = 16'h200;
			16'h42ed: y = 16'h200;
			16'h42ee: y = 16'h200;
			16'h42ef: y = 16'h200;
			16'h42f0: y = 16'h200;
			16'h42f1: y = 16'h200;
			16'h42f2: y = 16'h200;
			16'h42f3: y = 16'h200;
			16'h42f4: y = 16'h200;
			16'h42f5: y = 16'h200;
			16'h42f6: y = 16'h200;
			16'h42f7: y = 16'h200;
			16'h42f8: y = 16'h200;
			16'h42f9: y = 16'h200;
			16'h42fa: y = 16'h200;
			16'h42fb: y = 16'h200;
			16'h42fc: y = 16'h200;
			16'h42fd: y = 16'h200;
			16'h42fe: y = 16'h200;
			16'h42ff: y = 16'h200;
			16'h4300: y = 16'h200;
			16'h4301: y = 16'h200;
			16'h4302: y = 16'h200;
			16'h4303: y = 16'h200;
			16'h4304: y = 16'h200;
			16'h4305: y = 16'h200;
			16'h4306: y = 16'h200;
			16'h4307: y = 16'h200;
			16'h4308: y = 16'h200;
			16'h4309: y = 16'h200;
			16'h430a: y = 16'h200;
			16'h430b: y = 16'h200;
			16'h430c: y = 16'h200;
			16'h430d: y = 16'h200;
			16'h430e: y = 16'h200;
			16'h430f: y = 16'h200;
			16'h4310: y = 16'h200;
			16'h4311: y = 16'h200;
			16'h4312: y = 16'h200;
			16'h4313: y = 16'h200;
			16'h4314: y = 16'h200;
			16'h4315: y = 16'h200;
			16'h4316: y = 16'h200;
			16'h4317: y = 16'h200;
			16'h4318: y = 16'h200;
			16'h4319: y = 16'h200;
			16'h431a: y = 16'h200;
			16'h431b: y = 16'h200;
			16'h431c: y = 16'h200;
			16'h431d: y = 16'h200;
			16'h431e: y = 16'h200;
			16'h431f: y = 16'h200;
			16'h4320: y = 16'h200;
			16'h4321: y = 16'h200;
			16'h4322: y = 16'h200;
			16'h4323: y = 16'h200;
			16'h4324: y = 16'h200;
			16'h4325: y = 16'h200;
			16'h4326: y = 16'h200;
			16'h4327: y = 16'h200;
			16'h4328: y = 16'h200;
			16'h4329: y = 16'h200;
			16'h432a: y = 16'h200;
			16'h432b: y = 16'h200;
			16'h432c: y = 16'h200;
			16'h432d: y = 16'h200;
			16'h432e: y = 16'h200;
			16'h432f: y = 16'h200;
			16'h4330: y = 16'h200;
			16'h4331: y = 16'h200;
			16'h4332: y = 16'h200;
			16'h4333: y = 16'h200;
			16'h4334: y = 16'h200;
			16'h4335: y = 16'h200;
			16'h4336: y = 16'h200;
			16'h4337: y = 16'h200;
			16'h4338: y = 16'h200;
			16'h4339: y = 16'h200;
			16'h433a: y = 16'h200;
			16'h433b: y = 16'h200;
			16'h433c: y = 16'h200;
			16'h433d: y = 16'h200;
			16'h433e: y = 16'h200;
			16'h433f: y = 16'h200;
			16'h4340: y = 16'h200;
			16'h4341: y = 16'h200;
			16'h4342: y = 16'h200;
			16'h4343: y = 16'h200;
			16'h4344: y = 16'h200;
			16'h4345: y = 16'h200;
			16'h4346: y = 16'h200;
			16'h4347: y = 16'h200;
			16'h4348: y = 16'h200;
			16'h4349: y = 16'h200;
			16'h434a: y = 16'h200;
			16'h434b: y = 16'h200;
			16'h434c: y = 16'h200;
			16'h434d: y = 16'h200;
			16'h434e: y = 16'h200;
			16'h434f: y = 16'h200;
			16'h4350: y = 16'h200;
			16'h4351: y = 16'h200;
			16'h4352: y = 16'h200;
			16'h4353: y = 16'h200;
			16'h4354: y = 16'h200;
			16'h4355: y = 16'h200;
			16'h4356: y = 16'h200;
			16'h4357: y = 16'h200;
			16'h4358: y = 16'h200;
			16'h4359: y = 16'h200;
			16'h435a: y = 16'h200;
			16'h435b: y = 16'h200;
			16'h435c: y = 16'h200;
			16'h435d: y = 16'h200;
			16'h435e: y = 16'h200;
			16'h435f: y = 16'h200;
			16'h4360: y = 16'h200;
			16'h4361: y = 16'h200;
			16'h4362: y = 16'h200;
			16'h4363: y = 16'h200;
			16'h4364: y = 16'h200;
			16'h4365: y = 16'h200;
			16'h4366: y = 16'h200;
			16'h4367: y = 16'h200;
			16'h4368: y = 16'h200;
			16'h4369: y = 16'h200;
			16'h436a: y = 16'h200;
			16'h436b: y = 16'h200;
			16'h436c: y = 16'h200;
			16'h436d: y = 16'h200;
			16'h436e: y = 16'h200;
			16'h436f: y = 16'h200;
			16'h4370: y = 16'h200;
			16'h4371: y = 16'h200;
			16'h4372: y = 16'h200;
			16'h4373: y = 16'h200;
			16'h4374: y = 16'h200;
			16'h4375: y = 16'h200;
			16'h4376: y = 16'h200;
			16'h4377: y = 16'h200;
			16'h4378: y = 16'h200;
			16'h4379: y = 16'h200;
			16'h437a: y = 16'h200;
			16'h437b: y = 16'h200;
			16'h437c: y = 16'h200;
			16'h437d: y = 16'h200;
			16'h437e: y = 16'h200;
			16'h437f: y = 16'h200;
			16'h4380: y = 16'h200;
			16'h4381: y = 16'h200;
			16'h4382: y = 16'h200;
			16'h4383: y = 16'h200;
			16'h4384: y = 16'h200;
			16'h4385: y = 16'h200;
			16'h4386: y = 16'h200;
			16'h4387: y = 16'h200;
			16'h4388: y = 16'h200;
			16'h4389: y = 16'h200;
			16'h438a: y = 16'h200;
			16'h438b: y = 16'h200;
			16'h438c: y = 16'h200;
			16'h438d: y = 16'h200;
			16'h438e: y = 16'h200;
			16'h438f: y = 16'h200;
			16'h4390: y = 16'h200;
			16'h4391: y = 16'h200;
			16'h4392: y = 16'h200;
			16'h4393: y = 16'h200;
			16'h4394: y = 16'h200;
			16'h4395: y = 16'h200;
			16'h4396: y = 16'h200;
			16'h4397: y = 16'h200;
			16'h4398: y = 16'h200;
			16'h4399: y = 16'h200;
			16'h439a: y = 16'h200;
			16'h439b: y = 16'h200;
			16'h439c: y = 16'h200;
			16'h439d: y = 16'h200;
			16'h439e: y = 16'h200;
			16'h439f: y = 16'h200;
			16'h43a0: y = 16'h200;
			16'h43a1: y = 16'h200;
			16'h43a2: y = 16'h200;
			16'h43a3: y = 16'h200;
			16'h43a4: y = 16'h200;
			16'h43a5: y = 16'h200;
			16'h43a6: y = 16'h200;
			16'h43a7: y = 16'h200;
			16'h43a8: y = 16'h200;
			16'h43a9: y = 16'h200;
			16'h43aa: y = 16'h200;
			16'h43ab: y = 16'h200;
			16'h43ac: y = 16'h200;
			16'h43ad: y = 16'h200;
			16'h43ae: y = 16'h200;
			16'h43af: y = 16'h200;
			16'h43b0: y = 16'h200;
			16'h43b1: y = 16'h200;
			16'h43b2: y = 16'h200;
			16'h43b3: y = 16'h200;
			16'h43b4: y = 16'h200;
			16'h43b5: y = 16'h200;
			16'h43b6: y = 16'h200;
			16'h43b7: y = 16'h200;
			16'h43b8: y = 16'h200;
			16'h43b9: y = 16'h200;
			16'h43ba: y = 16'h200;
			16'h43bb: y = 16'h200;
			16'h43bc: y = 16'h200;
			16'h43bd: y = 16'h200;
			16'h43be: y = 16'h200;
			16'h43bf: y = 16'h200;
			16'h43c0: y = 16'h200;
			16'h43c1: y = 16'h200;
			16'h43c2: y = 16'h200;
			16'h43c3: y = 16'h200;
			16'h43c4: y = 16'h200;
			16'h43c5: y = 16'h200;
			16'h43c6: y = 16'h200;
			16'h43c7: y = 16'h200;
			16'h43c8: y = 16'h200;
			16'h43c9: y = 16'h200;
			16'h43ca: y = 16'h200;
			16'h43cb: y = 16'h200;
			16'h43cc: y = 16'h200;
			16'h43cd: y = 16'h200;
			16'h43ce: y = 16'h200;
			16'h43cf: y = 16'h200;
			16'h43d0: y = 16'h200;
			16'h43d1: y = 16'h200;
			16'h43d2: y = 16'h200;
			16'h43d3: y = 16'h200;
			16'h43d4: y = 16'h200;
			16'h43d5: y = 16'h200;
			16'h43d6: y = 16'h200;
			16'h43d7: y = 16'h200;
			16'h43d8: y = 16'h200;
			16'h43d9: y = 16'h200;
			16'h43da: y = 16'h200;
			16'h43db: y = 16'h200;
			16'h43dc: y = 16'h200;
			16'h43dd: y = 16'h200;
			16'h43de: y = 16'h200;
			16'h43df: y = 16'h200;
			16'h43e0: y = 16'h200;
			16'h43e1: y = 16'h200;
			16'h43e2: y = 16'h200;
			16'h43e3: y = 16'h200;
			16'h43e4: y = 16'h200;
			16'h43e5: y = 16'h200;
			16'h43e6: y = 16'h200;
			16'h43e7: y = 16'h200;
			16'h43e8: y = 16'h200;
			16'h43e9: y = 16'h200;
			16'h43ea: y = 16'h200;
			16'h43eb: y = 16'h200;
			16'h43ec: y = 16'h200;
			16'h43ed: y = 16'h200;
			16'h43ee: y = 16'h200;
			16'h43ef: y = 16'h200;
			16'h43f0: y = 16'h200;
			16'h43f1: y = 16'h200;
			16'h43f2: y = 16'h200;
			16'h43f3: y = 16'h200;
			16'h43f4: y = 16'h200;
			16'h43f5: y = 16'h200;
			16'h43f6: y = 16'h200;
			16'h43f7: y = 16'h200;
			16'h43f8: y = 16'h200;
			16'h43f9: y = 16'h200;
			16'h43fa: y = 16'h200;
			16'h43fb: y = 16'h200;
			16'h43fc: y = 16'h200;
			16'h43fd: y = 16'h200;
			16'h43fe: y = 16'h200;
			16'h43ff: y = 16'h200;
			16'h4400: y = 16'h200;
			16'h4401: y = 16'h200;
			16'h4402: y = 16'h200;
			16'h4403: y = 16'h200;
			16'h4404: y = 16'h200;
			16'h4405: y = 16'h200;
			16'h4406: y = 16'h200;
			16'h4407: y = 16'h200;
			16'h4408: y = 16'h200;
			16'h4409: y = 16'h200;
			16'h440a: y = 16'h200;
			16'h440b: y = 16'h200;
			16'h440c: y = 16'h200;
			16'h440d: y = 16'h200;
			16'h440e: y = 16'h200;
			16'h440f: y = 16'h200;
			16'h4410: y = 16'h200;
			16'h4411: y = 16'h200;
			16'h4412: y = 16'h200;
			16'h4413: y = 16'h200;
			16'h4414: y = 16'h200;
			16'h4415: y = 16'h200;
			16'h4416: y = 16'h200;
			16'h4417: y = 16'h200;
			16'h4418: y = 16'h200;
			16'h4419: y = 16'h200;
			16'h441a: y = 16'h200;
			16'h441b: y = 16'h200;
			16'h441c: y = 16'h200;
			16'h441d: y = 16'h200;
			16'h441e: y = 16'h200;
			16'h441f: y = 16'h200;
			16'h4420: y = 16'h200;
			16'h4421: y = 16'h200;
			16'h4422: y = 16'h200;
			16'h4423: y = 16'h200;
			16'h4424: y = 16'h200;
			16'h4425: y = 16'h200;
			16'h4426: y = 16'h200;
			16'h4427: y = 16'h200;
			16'h4428: y = 16'h200;
			16'h4429: y = 16'h200;
			16'h442a: y = 16'h200;
			16'h442b: y = 16'h200;
			16'h442c: y = 16'h200;
			16'h442d: y = 16'h200;
			16'h442e: y = 16'h200;
			16'h442f: y = 16'h200;
			16'h4430: y = 16'h200;
			16'h4431: y = 16'h200;
			16'h4432: y = 16'h200;
			16'h4433: y = 16'h200;
			16'h4434: y = 16'h200;
			16'h4435: y = 16'h200;
			16'h4436: y = 16'h200;
			16'h4437: y = 16'h200;
			16'h4438: y = 16'h200;
			16'h4439: y = 16'h200;
			16'h443a: y = 16'h200;
			16'h443b: y = 16'h200;
			16'h443c: y = 16'h200;
			16'h443d: y = 16'h200;
			16'h443e: y = 16'h200;
			16'h443f: y = 16'h200;
			16'h4440: y = 16'h200;
			16'h4441: y = 16'h200;
			16'h4442: y = 16'h200;
			16'h4443: y = 16'h200;
			16'h4444: y = 16'h200;
			16'h4445: y = 16'h200;
			16'h4446: y = 16'h200;
			16'h4447: y = 16'h200;
			16'h4448: y = 16'h200;
			16'h4449: y = 16'h200;
			16'h444a: y = 16'h200;
			16'h444b: y = 16'h200;
			16'h444c: y = 16'h200;
			16'h444d: y = 16'h200;
			16'h444e: y = 16'h200;
			16'h444f: y = 16'h200;
			16'h4450: y = 16'h200;
			16'h4451: y = 16'h200;
			16'h4452: y = 16'h200;
			16'h4453: y = 16'h200;
			16'h4454: y = 16'h200;
			16'h4455: y = 16'h200;
			16'h4456: y = 16'h200;
			16'h4457: y = 16'h200;
			16'h4458: y = 16'h200;
			16'h4459: y = 16'h200;
			16'h445a: y = 16'h200;
			16'h445b: y = 16'h200;
			16'h445c: y = 16'h200;
			16'h445d: y = 16'h200;
			16'h445e: y = 16'h200;
			16'h445f: y = 16'h200;
			16'h4460: y = 16'h200;
			16'h4461: y = 16'h200;
			16'h4462: y = 16'h200;
			16'h4463: y = 16'h200;
			16'h4464: y = 16'h200;
			16'h4465: y = 16'h200;
			16'h4466: y = 16'h200;
			16'h4467: y = 16'h200;
			16'h4468: y = 16'h200;
			16'h4469: y = 16'h200;
			16'h446a: y = 16'h200;
			16'h446b: y = 16'h200;
			16'h446c: y = 16'h200;
			16'h446d: y = 16'h200;
			16'h446e: y = 16'h200;
			16'h446f: y = 16'h200;
			16'h4470: y = 16'h200;
			16'h4471: y = 16'h200;
			16'h4472: y = 16'h200;
			16'h4473: y = 16'h200;
			16'h4474: y = 16'h200;
			16'h4475: y = 16'h200;
			16'h4476: y = 16'h200;
			16'h4477: y = 16'h200;
			16'h4478: y = 16'h200;
			16'h4479: y = 16'h200;
			16'h447a: y = 16'h200;
			16'h447b: y = 16'h200;
			16'h447c: y = 16'h200;
			16'h447d: y = 16'h200;
			16'h447e: y = 16'h200;
			16'h447f: y = 16'h200;
			16'h4480: y = 16'h200;
			16'h4481: y = 16'h200;
			16'h4482: y = 16'h200;
			16'h4483: y = 16'h200;
			16'h4484: y = 16'h200;
			16'h4485: y = 16'h200;
			16'h4486: y = 16'h200;
			16'h4487: y = 16'h200;
			16'h4488: y = 16'h200;
			16'h4489: y = 16'h200;
			16'h448a: y = 16'h200;
			16'h448b: y = 16'h200;
			16'h448c: y = 16'h200;
			16'h448d: y = 16'h200;
			16'h448e: y = 16'h200;
			16'h448f: y = 16'h200;
			16'h4490: y = 16'h200;
			16'h4491: y = 16'h200;
			16'h4492: y = 16'h200;
			16'h4493: y = 16'h200;
			16'h4494: y = 16'h200;
			16'h4495: y = 16'h200;
			16'h4496: y = 16'h200;
			16'h4497: y = 16'h200;
			16'h4498: y = 16'h200;
			16'h4499: y = 16'h200;
			16'h449a: y = 16'h200;
			16'h449b: y = 16'h200;
			16'h449c: y = 16'h200;
			16'h449d: y = 16'h200;
			16'h449e: y = 16'h200;
			16'h449f: y = 16'h200;
			16'h44a0: y = 16'h200;
			16'h44a1: y = 16'h200;
			16'h44a2: y = 16'h200;
			16'h44a3: y = 16'h200;
			16'h44a4: y = 16'h200;
			16'h44a5: y = 16'h200;
			16'h44a6: y = 16'h200;
			16'h44a7: y = 16'h200;
			16'h44a8: y = 16'h200;
			16'h44a9: y = 16'h200;
			16'h44aa: y = 16'h200;
			16'h44ab: y = 16'h200;
			16'h44ac: y = 16'h200;
			16'h44ad: y = 16'h200;
			16'h44ae: y = 16'h200;
			16'h44af: y = 16'h200;
			16'h44b0: y = 16'h200;
			16'h44b1: y = 16'h200;
			16'h44b2: y = 16'h200;
			16'h44b3: y = 16'h200;
			16'h44b4: y = 16'h200;
			16'h44b5: y = 16'h200;
			16'h44b6: y = 16'h200;
			16'h44b7: y = 16'h200;
			16'h44b8: y = 16'h200;
			16'h44b9: y = 16'h200;
			16'h44ba: y = 16'h200;
			16'h44bb: y = 16'h200;
			16'h44bc: y = 16'h200;
			16'h44bd: y = 16'h200;
			16'h44be: y = 16'h200;
			16'h44bf: y = 16'h200;
			16'h44c0: y = 16'h200;
			16'h44c1: y = 16'h200;
			16'h44c2: y = 16'h200;
			16'h44c3: y = 16'h200;
			16'h44c4: y = 16'h200;
			16'h44c5: y = 16'h200;
			16'h44c6: y = 16'h200;
			16'h44c7: y = 16'h200;
			16'h44c8: y = 16'h200;
			16'h44c9: y = 16'h200;
			16'h44ca: y = 16'h200;
			16'h44cb: y = 16'h200;
			16'h44cc: y = 16'h200;
			16'h44cd: y = 16'h200;
			16'h44ce: y = 16'h200;
			16'h44cf: y = 16'h200;
			16'h44d0: y = 16'h200;
			16'h44d1: y = 16'h200;
			16'h44d2: y = 16'h200;
			16'h44d3: y = 16'h200;
			16'h44d4: y = 16'h200;
			16'h44d5: y = 16'h200;
			16'h44d6: y = 16'h200;
			16'h44d7: y = 16'h200;
			16'h44d8: y = 16'h200;
			16'h44d9: y = 16'h200;
			16'h44da: y = 16'h200;
			16'h44db: y = 16'h200;
			16'h44dc: y = 16'h200;
			16'h44dd: y = 16'h200;
			16'h44de: y = 16'h200;
			16'h44df: y = 16'h200;
			16'h44e0: y = 16'h200;
			16'h44e1: y = 16'h200;
			16'h44e2: y = 16'h200;
			16'h44e3: y = 16'h200;
			16'h44e4: y = 16'h200;
			16'h44e5: y = 16'h200;
			16'h44e6: y = 16'h200;
			16'h44e7: y = 16'h200;
			16'h44e8: y = 16'h200;
			16'h44e9: y = 16'h200;
			16'h44ea: y = 16'h200;
			16'h44eb: y = 16'h200;
			16'h44ec: y = 16'h200;
			16'h44ed: y = 16'h200;
			16'h44ee: y = 16'h200;
			16'h44ef: y = 16'h200;
			16'h44f0: y = 16'h200;
			16'h44f1: y = 16'h200;
			16'h44f2: y = 16'h200;
			16'h44f3: y = 16'h200;
			16'h44f4: y = 16'h200;
			16'h44f5: y = 16'h200;
			16'h44f6: y = 16'h200;
			16'h44f7: y = 16'h200;
			16'h44f8: y = 16'h200;
			16'h44f9: y = 16'h200;
			16'h44fa: y = 16'h200;
			16'h44fb: y = 16'h200;
			16'h44fc: y = 16'h200;
			16'h44fd: y = 16'h200;
			16'h44fe: y = 16'h200;
			16'h44ff: y = 16'h200;
			16'h4500: y = 16'h200;
			16'h4501: y = 16'h200;
			16'h4502: y = 16'h200;
			16'h4503: y = 16'h200;
			16'h4504: y = 16'h200;
			16'h4505: y = 16'h200;
			16'h4506: y = 16'h200;
			16'h4507: y = 16'h200;
			16'h4508: y = 16'h200;
			16'h4509: y = 16'h200;
			16'h450a: y = 16'h200;
			16'h450b: y = 16'h200;
			16'h450c: y = 16'h200;
			16'h450d: y = 16'h200;
			16'h450e: y = 16'h200;
			16'h450f: y = 16'h200;
			16'h4510: y = 16'h200;
			16'h4511: y = 16'h200;
			16'h4512: y = 16'h200;
			16'h4513: y = 16'h200;
			16'h4514: y = 16'h200;
			16'h4515: y = 16'h200;
			16'h4516: y = 16'h200;
			16'h4517: y = 16'h200;
			16'h4518: y = 16'h200;
			16'h4519: y = 16'h200;
			16'h451a: y = 16'h200;
			16'h451b: y = 16'h200;
			16'h451c: y = 16'h200;
			16'h451d: y = 16'h200;
			16'h451e: y = 16'h200;
			16'h451f: y = 16'h200;
			16'h4520: y = 16'h200;
			16'h4521: y = 16'h200;
			16'h4522: y = 16'h200;
			16'h4523: y = 16'h200;
			16'h4524: y = 16'h200;
			16'h4525: y = 16'h200;
			16'h4526: y = 16'h200;
			16'h4527: y = 16'h200;
			16'h4528: y = 16'h200;
			16'h4529: y = 16'h200;
			16'h452a: y = 16'h200;
			16'h452b: y = 16'h200;
			16'h452c: y = 16'h200;
			16'h452d: y = 16'h200;
			16'h452e: y = 16'h200;
			16'h452f: y = 16'h200;
			16'h4530: y = 16'h200;
			16'h4531: y = 16'h200;
			16'h4532: y = 16'h200;
			16'h4533: y = 16'h200;
			16'h4534: y = 16'h200;
			16'h4535: y = 16'h200;
			16'h4536: y = 16'h200;
			16'h4537: y = 16'h200;
			16'h4538: y = 16'h200;
			16'h4539: y = 16'h200;
			16'h453a: y = 16'h200;
			16'h453b: y = 16'h200;
			16'h453c: y = 16'h200;
			16'h453d: y = 16'h200;
			16'h453e: y = 16'h200;
			16'h453f: y = 16'h200;
			16'h4540: y = 16'h200;
			16'h4541: y = 16'h200;
			16'h4542: y = 16'h200;
			16'h4543: y = 16'h200;
			16'h4544: y = 16'h200;
			16'h4545: y = 16'h200;
			16'h4546: y = 16'h200;
			16'h4547: y = 16'h200;
			16'h4548: y = 16'h200;
			16'h4549: y = 16'h200;
			16'h454a: y = 16'h200;
			16'h454b: y = 16'h200;
			16'h454c: y = 16'h200;
			16'h454d: y = 16'h200;
			16'h454e: y = 16'h200;
			16'h454f: y = 16'h200;
			16'h4550: y = 16'h200;
			16'h4551: y = 16'h200;
			16'h4552: y = 16'h200;
			16'h4553: y = 16'h200;
			16'h4554: y = 16'h200;
			16'h4555: y = 16'h200;
			16'h4556: y = 16'h200;
			16'h4557: y = 16'h200;
			16'h4558: y = 16'h200;
			16'h4559: y = 16'h200;
			16'h455a: y = 16'h200;
			16'h455b: y = 16'h200;
			16'h455c: y = 16'h200;
			16'h455d: y = 16'h200;
			16'h455e: y = 16'h200;
			16'h455f: y = 16'h200;
			16'h4560: y = 16'h200;
			16'h4561: y = 16'h200;
			16'h4562: y = 16'h200;
			16'h4563: y = 16'h200;
			16'h4564: y = 16'h200;
			16'h4565: y = 16'h200;
			16'h4566: y = 16'h200;
			16'h4567: y = 16'h200;
			16'h4568: y = 16'h200;
			16'h4569: y = 16'h200;
			16'h456a: y = 16'h200;
			16'h456b: y = 16'h200;
			16'h456c: y = 16'h200;
			16'h456d: y = 16'h200;
			16'h456e: y = 16'h200;
			16'h456f: y = 16'h200;
			16'h4570: y = 16'h200;
			16'h4571: y = 16'h200;
			16'h4572: y = 16'h200;
			16'h4573: y = 16'h200;
			16'h4574: y = 16'h200;
			16'h4575: y = 16'h200;
			16'h4576: y = 16'h200;
			16'h4577: y = 16'h200;
			16'h4578: y = 16'h200;
			16'h4579: y = 16'h200;
			16'h457a: y = 16'h200;
			16'h457b: y = 16'h200;
			16'h457c: y = 16'h200;
			16'h457d: y = 16'h200;
			16'h457e: y = 16'h200;
			16'h457f: y = 16'h200;
			16'h4580: y = 16'h200;
			16'h4581: y = 16'h200;
			16'h4582: y = 16'h200;
			16'h4583: y = 16'h200;
			16'h4584: y = 16'h200;
			16'h4585: y = 16'h200;
			16'h4586: y = 16'h200;
			16'h4587: y = 16'h200;
			16'h4588: y = 16'h200;
			16'h4589: y = 16'h200;
			16'h458a: y = 16'h200;
			16'h458b: y = 16'h200;
			16'h458c: y = 16'h200;
			16'h458d: y = 16'h200;
			16'h458e: y = 16'h200;
			16'h458f: y = 16'h200;
			16'h4590: y = 16'h200;
			16'h4591: y = 16'h200;
			16'h4592: y = 16'h200;
			16'h4593: y = 16'h200;
			16'h4594: y = 16'h200;
			16'h4595: y = 16'h200;
			16'h4596: y = 16'h200;
			16'h4597: y = 16'h200;
			16'h4598: y = 16'h200;
			16'h4599: y = 16'h200;
			16'h459a: y = 16'h200;
			16'h459b: y = 16'h200;
			16'h459c: y = 16'h200;
			16'h459d: y = 16'h200;
			16'h459e: y = 16'h200;
			16'h459f: y = 16'h200;
			16'h45a0: y = 16'h200;
			16'h45a1: y = 16'h200;
			16'h45a2: y = 16'h200;
			16'h45a3: y = 16'h200;
			16'h45a4: y = 16'h200;
			16'h45a5: y = 16'h200;
			16'h45a6: y = 16'h200;
			16'h45a7: y = 16'h200;
			16'h45a8: y = 16'h200;
			16'h45a9: y = 16'h200;
			16'h45aa: y = 16'h200;
			16'h45ab: y = 16'h200;
			16'h45ac: y = 16'h200;
			16'h45ad: y = 16'h200;
			16'h45ae: y = 16'h200;
			16'h45af: y = 16'h200;
			16'h45b0: y = 16'h200;
			16'h45b1: y = 16'h200;
			16'h45b2: y = 16'h200;
			16'h45b3: y = 16'h200;
			16'h45b4: y = 16'h200;
			16'h45b5: y = 16'h200;
			16'h45b6: y = 16'h200;
			16'h45b7: y = 16'h200;
			16'h45b8: y = 16'h200;
			16'h45b9: y = 16'h200;
			16'h45ba: y = 16'h200;
			16'h45bb: y = 16'h200;
			16'h45bc: y = 16'h200;
			16'h45bd: y = 16'h200;
			16'h45be: y = 16'h200;
			16'h45bf: y = 16'h200;
			16'h45c0: y = 16'h200;
			16'h45c1: y = 16'h200;
			16'h45c2: y = 16'h200;
			16'h45c3: y = 16'h200;
			16'h45c4: y = 16'h200;
			16'h45c5: y = 16'h200;
			16'h45c6: y = 16'h200;
			16'h45c7: y = 16'h200;
			16'h45c8: y = 16'h200;
			16'h45c9: y = 16'h200;
			16'h45ca: y = 16'h200;
			16'h45cb: y = 16'h200;
			16'h45cc: y = 16'h200;
			16'h45cd: y = 16'h200;
			16'h45ce: y = 16'h200;
			16'h45cf: y = 16'h200;
			16'h45d0: y = 16'h200;
			16'h45d1: y = 16'h200;
			16'h45d2: y = 16'h200;
			16'h45d3: y = 16'h200;
			16'h45d4: y = 16'h200;
			16'h45d5: y = 16'h200;
			16'h45d6: y = 16'h200;
			16'h45d7: y = 16'h200;
			16'h45d8: y = 16'h200;
			16'h45d9: y = 16'h200;
			16'h45da: y = 16'h200;
			16'h45db: y = 16'h200;
			16'h45dc: y = 16'h200;
			16'h45dd: y = 16'h200;
			16'h45de: y = 16'h200;
			16'h45df: y = 16'h200;
			16'h45e0: y = 16'h200;
			16'h45e1: y = 16'h200;
			16'h45e2: y = 16'h200;
			16'h45e3: y = 16'h200;
			16'h45e4: y = 16'h200;
			16'h45e5: y = 16'h200;
			16'h45e6: y = 16'h200;
			16'h45e7: y = 16'h200;
			16'h45e8: y = 16'h200;
			16'h45e9: y = 16'h200;
			16'h45ea: y = 16'h200;
			16'h45eb: y = 16'h200;
			16'h45ec: y = 16'h200;
			16'h45ed: y = 16'h200;
			16'h45ee: y = 16'h200;
			16'h45ef: y = 16'h200;
			16'h45f0: y = 16'h200;
			16'h45f1: y = 16'h200;
			16'h45f2: y = 16'h200;
			16'h45f3: y = 16'h200;
			16'h45f4: y = 16'h200;
			16'h45f5: y = 16'h200;
			16'h45f6: y = 16'h200;
			16'h45f7: y = 16'h200;
			16'h45f8: y = 16'h200;
			16'h45f9: y = 16'h200;
			16'h45fa: y = 16'h200;
			16'h45fb: y = 16'h200;
			16'h45fc: y = 16'h200;
			16'h45fd: y = 16'h200;
			16'h45fe: y = 16'h200;
			16'h45ff: y = 16'h200;
			16'h4600: y = 16'h200;
			16'h4601: y = 16'h200;
			16'h4602: y = 16'h200;
			16'h4603: y = 16'h200;
			16'h4604: y = 16'h200;
			16'h4605: y = 16'h200;
			16'h4606: y = 16'h200;
			16'h4607: y = 16'h200;
			16'h4608: y = 16'h200;
			16'h4609: y = 16'h200;
			16'h460a: y = 16'h200;
			16'h460b: y = 16'h200;
			16'h460c: y = 16'h200;
			16'h460d: y = 16'h200;
			16'h460e: y = 16'h200;
			16'h460f: y = 16'h200;
			16'h4610: y = 16'h200;
			16'h4611: y = 16'h200;
			16'h4612: y = 16'h200;
			16'h4613: y = 16'h200;
			16'h4614: y = 16'h200;
			16'h4615: y = 16'h200;
			16'h4616: y = 16'h200;
			16'h4617: y = 16'h200;
			16'h4618: y = 16'h200;
			16'h4619: y = 16'h200;
			16'h461a: y = 16'h200;
			16'h461b: y = 16'h200;
			16'h461c: y = 16'h200;
			16'h461d: y = 16'h200;
			16'h461e: y = 16'h200;
			16'h461f: y = 16'h200;
			16'h4620: y = 16'h200;
			16'h4621: y = 16'h200;
			16'h4622: y = 16'h200;
			16'h4623: y = 16'h200;
			16'h4624: y = 16'h200;
			16'h4625: y = 16'h200;
			16'h4626: y = 16'h200;
			16'h4627: y = 16'h200;
			16'h4628: y = 16'h200;
			16'h4629: y = 16'h200;
			16'h462a: y = 16'h200;
			16'h462b: y = 16'h200;
			16'h462c: y = 16'h200;
			16'h462d: y = 16'h200;
			16'h462e: y = 16'h200;
			16'h462f: y = 16'h200;
			16'h4630: y = 16'h200;
			16'h4631: y = 16'h200;
			16'h4632: y = 16'h200;
			16'h4633: y = 16'h200;
			16'h4634: y = 16'h200;
			16'h4635: y = 16'h200;
			16'h4636: y = 16'h200;
			16'h4637: y = 16'h200;
			16'h4638: y = 16'h200;
			16'h4639: y = 16'h200;
			16'h463a: y = 16'h200;
			16'h463b: y = 16'h200;
			16'h463c: y = 16'h200;
			16'h463d: y = 16'h200;
			16'h463e: y = 16'h200;
			16'h463f: y = 16'h200;
			16'h4640: y = 16'h200;
			16'h4641: y = 16'h200;
			16'h4642: y = 16'h200;
			16'h4643: y = 16'h200;
			16'h4644: y = 16'h200;
			16'h4645: y = 16'h200;
			16'h4646: y = 16'h200;
			16'h4647: y = 16'h200;
			16'h4648: y = 16'h200;
			16'h4649: y = 16'h200;
			16'h464a: y = 16'h200;
			16'h464b: y = 16'h200;
			16'h464c: y = 16'h200;
			16'h464d: y = 16'h200;
			16'h464e: y = 16'h200;
			16'h464f: y = 16'h200;
			16'h4650: y = 16'h200;
			16'h4651: y = 16'h200;
			16'h4652: y = 16'h200;
			16'h4653: y = 16'h200;
			16'h4654: y = 16'h200;
			16'h4655: y = 16'h200;
			16'h4656: y = 16'h200;
			16'h4657: y = 16'h200;
			16'h4658: y = 16'h200;
			16'h4659: y = 16'h200;
			16'h465a: y = 16'h200;
			16'h465b: y = 16'h200;
			16'h465c: y = 16'h200;
			16'h465d: y = 16'h200;
			16'h465e: y = 16'h200;
			16'h465f: y = 16'h200;
			16'h4660: y = 16'h200;
			16'h4661: y = 16'h200;
			16'h4662: y = 16'h200;
			16'h4663: y = 16'h200;
			16'h4664: y = 16'h200;
			16'h4665: y = 16'h200;
			16'h4666: y = 16'h200;
			16'h4667: y = 16'h200;
			16'h4668: y = 16'h200;
			16'h4669: y = 16'h200;
			16'h466a: y = 16'h200;
			16'h466b: y = 16'h200;
			16'h466c: y = 16'h200;
			16'h466d: y = 16'h200;
			16'h466e: y = 16'h200;
			16'h466f: y = 16'h200;
			16'h4670: y = 16'h200;
			16'h4671: y = 16'h200;
			16'h4672: y = 16'h200;
			16'h4673: y = 16'h200;
			16'h4674: y = 16'h200;
			16'h4675: y = 16'h200;
			16'h4676: y = 16'h200;
			16'h4677: y = 16'h200;
			16'h4678: y = 16'h200;
			16'h4679: y = 16'h200;
			16'h467a: y = 16'h200;
			16'h467b: y = 16'h200;
			16'h467c: y = 16'h200;
			16'h467d: y = 16'h200;
			16'h467e: y = 16'h200;
			16'h467f: y = 16'h200;
			16'h4680: y = 16'h200;
			16'h4681: y = 16'h200;
			16'h4682: y = 16'h200;
			16'h4683: y = 16'h200;
			16'h4684: y = 16'h200;
			16'h4685: y = 16'h200;
			16'h4686: y = 16'h200;
			16'h4687: y = 16'h200;
			16'h4688: y = 16'h200;
			16'h4689: y = 16'h200;
			16'h468a: y = 16'h200;
			16'h468b: y = 16'h200;
			16'h468c: y = 16'h200;
			16'h468d: y = 16'h200;
			16'h468e: y = 16'h200;
			16'h468f: y = 16'h200;
			16'h4690: y = 16'h200;
			16'h4691: y = 16'h200;
			16'h4692: y = 16'h200;
			16'h4693: y = 16'h200;
			16'h4694: y = 16'h200;
			16'h4695: y = 16'h200;
			16'h4696: y = 16'h200;
			16'h4697: y = 16'h200;
			16'h4698: y = 16'h200;
			16'h4699: y = 16'h200;
			16'h469a: y = 16'h200;
			16'h469b: y = 16'h200;
			16'h469c: y = 16'h200;
			16'h469d: y = 16'h200;
			16'h469e: y = 16'h200;
			16'h469f: y = 16'h200;
			16'h46a0: y = 16'h200;
			16'h46a1: y = 16'h200;
			16'h46a2: y = 16'h200;
			16'h46a3: y = 16'h200;
			16'h46a4: y = 16'h200;
			16'h46a5: y = 16'h200;
			16'h46a6: y = 16'h200;
			16'h46a7: y = 16'h200;
			16'h46a8: y = 16'h200;
			16'h46a9: y = 16'h200;
			16'h46aa: y = 16'h200;
			16'h46ab: y = 16'h200;
			16'h46ac: y = 16'h200;
			16'h46ad: y = 16'h200;
			16'h46ae: y = 16'h200;
			16'h46af: y = 16'h200;
			16'h46b0: y = 16'h200;
			16'h46b1: y = 16'h200;
			16'h46b2: y = 16'h200;
			16'h46b3: y = 16'h200;
			16'h46b4: y = 16'h200;
			16'h46b5: y = 16'h200;
			16'h46b6: y = 16'h200;
			16'h46b7: y = 16'h200;
			16'h46b8: y = 16'h200;
			16'h46b9: y = 16'h200;
			16'h46ba: y = 16'h200;
			16'h46bb: y = 16'h200;
			16'h46bc: y = 16'h200;
			16'h46bd: y = 16'h200;
			16'h46be: y = 16'h200;
			16'h46bf: y = 16'h200;
			16'h46c0: y = 16'h200;
			16'h46c1: y = 16'h200;
			16'h46c2: y = 16'h200;
			16'h46c3: y = 16'h200;
			16'h46c4: y = 16'h200;
			16'h46c5: y = 16'h200;
			16'h46c6: y = 16'h200;
			16'h46c7: y = 16'h200;
			16'h46c8: y = 16'h200;
			16'h46c9: y = 16'h200;
			16'h46ca: y = 16'h200;
			16'h46cb: y = 16'h200;
			16'h46cc: y = 16'h200;
			16'h46cd: y = 16'h200;
			16'h46ce: y = 16'h200;
			16'h46cf: y = 16'h200;
			16'h46d0: y = 16'h200;
			16'h46d1: y = 16'h200;
			16'h46d2: y = 16'h200;
			16'h46d3: y = 16'h200;
			16'h46d4: y = 16'h200;
			16'h46d5: y = 16'h200;
			16'h46d6: y = 16'h200;
			16'h46d7: y = 16'h200;
			16'h46d8: y = 16'h200;
			16'h46d9: y = 16'h200;
			16'h46da: y = 16'h200;
			16'h46db: y = 16'h200;
			16'h46dc: y = 16'h200;
			16'h46dd: y = 16'h200;
			16'h46de: y = 16'h200;
			16'h46df: y = 16'h200;
			16'h46e0: y = 16'h200;
			16'h46e1: y = 16'h200;
			16'h46e2: y = 16'h200;
			16'h46e3: y = 16'h200;
			16'h46e4: y = 16'h200;
			16'h46e5: y = 16'h200;
			16'h46e6: y = 16'h200;
			16'h46e7: y = 16'h200;
			16'h46e8: y = 16'h200;
			16'h46e9: y = 16'h200;
			16'h46ea: y = 16'h200;
			16'h46eb: y = 16'h200;
			16'h46ec: y = 16'h200;
			16'h46ed: y = 16'h200;
			16'h46ee: y = 16'h200;
			16'h46ef: y = 16'h200;
			16'h46f0: y = 16'h200;
			16'h46f1: y = 16'h200;
			16'h46f2: y = 16'h200;
			16'h46f3: y = 16'h200;
			16'h46f4: y = 16'h200;
			16'h46f5: y = 16'h200;
			16'h46f6: y = 16'h200;
			16'h46f7: y = 16'h200;
			16'h46f8: y = 16'h200;
			16'h46f9: y = 16'h200;
			16'h46fa: y = 16'h200;
			16'h46fb: y = 16'h200;
			16'h46fc: y = 16'h200;
			16'h46fd: y = 16'h200;
			16'h46fe: y = 16'h200;
			16'h46ff: y = 16'h200;
			16'h4700: y = 16'h200;
			16'h4701: y = 16'h200;
			16'h4702: y = 16'h200;
			16'h4703: y = 16'h200;
			16'h4704: y = 16'h200;
			16'h4705: y = 16'h200;
			16'h4706: y = 16'h200;
			16'h4707: y = 16'h200;
			16'h4708: y = 16'h200;
			16'h4709: y = 16'h200;
			16'h470a: y = 16'h200;
			16'h470b: y = 16'h200;
			16'h470c: y = 16'h200;
			16'h470d: y = 16'h200;
			16'h470e: y = 16'h200;
			16'h470f: y = 16'h200;
			16'h4710: y = 16'h200;
			16'h4711: y = 16'h200;
			16'h4712: y = 16'h200;
			16'h4713: y = 16'h200;
			16'h4714: y = 16'h200;
			16'h4715: y = 16'h200;
			16'h4716: y = 16'h200;
			16'h4717: y = 16'h200;
			16'h4718: y = 16'h200;
			16'h4719: y = 16'h200;
			16'h471a: y = 16'h200;
			16'h471b: y = 16'h200;
			16'h471c: y = 16'h200;
			16'h471d: y = 16'h200;
			16'h471e: y = 16'h200;
			16'h471f: y = 16'h200;
			16'h4720: y = 16'h200;
			16'h4721: y = 16'h200;
			16'h4722: y = 16'h200;
			16'h4723: y = 16'h200;
			16'h4724: y = 16'h200;
			16'h4725: y = 16'h200;
			16'h4726: y = 16'h200;
			16'h4727: y = 16'h200;
			16'h4728: y = 16'h200;
			16'h4729: y = 16'h200;
			16'h472a: y = 16'h200;
			16'h472b: y = 16'h200;
			16'h472c: y = 16'h200;
			16'h472d: y = 16'h200;
			16'h472e: y = 16'h200;
			16'h472f: y = 16'h200;
			16'h4730: y = 16'h200;
			16'h4731: y = 16'h200;
			16'h4732: y = 16'h200;
			16'h4733: y = 16'h200;
			16'h4734: y = 16'h200;
			16'h4735: y = 16'h200;
			16'h4736: y = 16'h200;
			16'h4737: y = 16'h200;
			16'h4738: y = 16'h200;
			16'h4739: y = 16'h200;
			16'h473a: y = 16'h200;
			16'h473b: y = 16'h200;
			16'h473c: y = 16'h200;
			16'h473d: y = 16'h200;
			16'h473e: y = 16'h200;
			16'h473f: y = 16'h200;
			16'h4740: y = 16'h200;
			16'h4741: y = 16'h200;
			16'h4742: y = 16'h200;
			16'h4743: y = 16'h200;
			16'h4744: y = 16'h200;
			16'h4745: y = 16'h200;
			16'h4746: y = 16'h200;
			16'h4747: y = 16'h200;
			16'h4748: y = 16'h200;
			16'h4749: y = 16'h200;
			16'h474a: y = 16'h200;
			16'h474b: y = 16'h200;
			16'h474c: y = 16'h200;
			16'h474d: y = 16'h200;
			16'h474e: y = 16'h200;
			16'h474f: y = 16'h200;
			16'h4750: y = 16'h200;
			16'h4751: y = 16'h200;
			16'h4752: y = 16'h200;
			16'h4753: y = 16'h200;
			16'h4754: y = 16'h200;
			16'h4755: y = 16'h200;
			16'h4756: y = 16'h200;
			16'h4757: y = 16'h200;
			16'h4758: y = 16'h200;
			16'h4759: y = 16'h200;
			16'h475a: y = 16'h200;
			16'h475b: y = 16'h200;
			16'h475c: y = 16'h200;
			16'h475d: y = 16'h200;
			16'h475e: y = 16'h200;
			16'h475f: y = 16'h200;
			16'h4760: y = 16'h200;
			16'h4761: y = 16'h200;
			16'h4762: y = 16'h200;
			16'h4763: y = 16'h200;
			16'h4764: y = 16'h200;
			16'h4765: y = 16'h200;
			16'h4766: y = 16'h200;
			16'h4767: y = 16'h200;
			16'h4768: y = 16'h200;
			16'h4769: y = 16'h200;
			16'h476a: y = 16'h200;
			16'h476b: y = 16'h200;
			16'h476c: y = 16'h200;
			16'h476d: y = 16'h200;
			16'h476e: y = 16'h200;
			16'h476f: y = 16'h200;
			16'h4770: y = 16'h200;
			16'h4771: y = 16'h200;
			16'h4772: y = 16'h200;
			16'h4773: y = 16'h200;
			16'h4774: y = 16'h200;
			16'h4775: y = 16'h200;
			16'h4776: y = 16'h200;
			16'h4777: y = 16'h200;
			16'h4778: y = 16'h200;
			16'h4779: y = 16'h200;
			16'h477a: y = 16'h200;
			16'h477b: y = 16'h200;
			16'h477c: y = 16'h200;
			16'h477d: y = 16'h200;
			16'h477e: y = 16'h200;
			16'h477f: y = 16'h200;
			16'h4780: y = 16'h200;
			16'h4781: y = 16'h200;
			16'h4782: y = 16'h200;
			16'h4783: y = 16'h200;
			16'h4784: y = 16'h200;
			16'h4785: y = 16'h200;
			16'h4786: y = 16'h200;
			16'h4787: y = 16'h200;
			16'h4788: y = 16'h200;
			16'h4789: y = 16'h200;
			16'h478a: y = 16'h200;
			16'h478b: y = 16'h200;
			16'h478c: y = 16'h200;
			16'h478d: y = 16'h200;
			16'h478e: y = 16'h200;
			16'h478f: y = 16'h200;
			16'h4790: y = 16'h200;
			16'h4791: y = 16'h200;
			16'h4792: y = 16'h200;
			16'h4793: y = 16'h200;
			16'h4794: y = 16'h200;
			16'h4795: y = 16'h200;
			16'h4796: y = 16'h200;
			16'h4797: y = 16'h200;
			16'h4798: y = 16'h200;
			16'h4799: y = 16'h200;
			16'h479a: y = 16'h200;
			16'h479b: y = 16'h200;
			16'h479c: y = 16'h200;
			16'h479d: y = 16'h200;
			16'h479e: y = 16'h200;
			16'h479f: y = 16'h200;
			16'h47a0: y = 16'h200;
			16'h47a1: y = 16'h200;
			16'h47a2: y = 16'h200;
			16'h47a3: y = 16'h200;
			16'h47a4: y = 16'h200;
			16'h47a5: y = 16'h200;
			16'h47a6: y = 16'h200;
			16'h47a7: y = 16'h200;
			16'h47a8: y = 16'h200;
			16'h47a9: y = 16'h200;
			16'h47aa: y = 16'h200;
			16'h47ab: y = 16'h200;
			16'h47ac: y = 16'h200;
			16'h47ad: y = 16'h200;
			16'h47ae: y = 16'h200;
			16'h47af: y = 16'h200;
			16'h47b0: y = 16'h200;
			16'h47b1: y = 16'h200;
			16'h47b2: y = 16'h200;
			16'h47b3: y = 16'h200;
			16'h47b4: y = 16'h200;
			16'h47b5: y = 16'h200;
			16'h47b6: y = 16'h200;
			16'h47b7: y = 16'h200;
			16'h47b8: y = 16'h200;
			16'h47b9: y = 16'h200;
			16'h47ba: y = 16'h200;
			16'h47bb: y = 16'h200;
			16'h47bc: y = 16'h200;
			16'h47bd: y = 16'h200;
			16'h47be: y = 16'h200;
			16'h47bf: y = 16'h200;
			16'h47c0: y = 16'h200;
			16'h47c1: y = 16'h200;
			16'h47c2: y = 16'h200;
			16'h47c3: y = 16'h200;
			16'h47c4: y = 16'h200;
			16'h47c5: y = 16'h200;
			16'h47c6: y = 16'h200;
			16'h47c7: y = 16'h200;
			16'h47c8: y = 16'h200;
			16'h47c9: y = 16'h200;
			16'h47ca: y = 16'h200;
			16'h47cb: y = 16'h200;
			16'h47cc: y = 16'h200;
			16'h47cd: y = 16'h200;
			16'h47ce: y = 16'h200;
			16'h47cf: y = 16'h200;
			16'h47d0: y = 16'h200;
			16'h47d1: y = 16'h200;
			16'h47d2: y = 16'h200;
			16'h47d3: y = 16'h200;
			16'h47d4: y = 16'h200;
			16'h47d5: y = 16'h200;
			16'h47d6: y = 16'h200;
			16'h47d7: y = 16'h200;
			16'h47d8: y = 16'h200;
			16'h47d9: y = 16'h200;
			16'h47da: y = 16'h200;
			16'h47db: y = 16'h200;
			16'h47dc: y = 16'h200;
			16'h47dd: y = 16'h200;
			16'h47de: y = 16'h200;
			16'h47df: y = 16'h200;
			16'h47e0: y = 16'h200;
			16'h47e1: y = 16'h200;
			16'h47e2: y = 16'h200;
			16'h47e3: y = 16'h200;
			16'h47e4: y = 16'h200;
			16'h47e5: y = 16'h200;
			16'h47e6: y = 16'h200;
			16'h47e7: y = 16'h200;
			16'h47e8: y = 16'h200;
			16'h47e9: y = 16'h200;
			16'h47ea: y = 16'h200;
			16'h47eb: y = 16'h200;
			16'h47ec: y = 16'h200;
			16'h47ed: y = 16'h200;
			16'h47ee: y = 16'h200;
			16'h47ef: y = 16'h200;
			16'h47f0: y = 16'h200;
			16'h47f1: y = 16'h200;
			16'h47f2: y = 16'h200;
			16'h47f3: y = 16'h200;
			16'h47f4: y = 16'h200;
			16'h47f5: y = 16'h200;
			16'h47f6: y = 16'h200;
			16'h47f7: y = 16'h200;
			16'h47f8: y = 16'h200;
			16'h47f9: y = 16'h200;
			16'h47fa: y = 16'h200;
			16'h47fb: y = 16'h200;
			16'h47fc: y = 16'h200;
			16'h47fd: y = 16'h200;
			16'h47fe: y = 16'h200;
			16'h47ff: y = 16'h200;
			16'h4800: y = 16'h200;
			16'h4801: y = 16'h200;
			16'h4802: y = 16'h200;
			16'h4803: y = 16'h200;
			16'h4804: y = 16'h200;
			16'h4805: y = 16'h200;
			16'h4806: y = 16'h200;
			16'h4807: y = 16'h200;
			16'h4808: y = 16'h200;
			16'h4809: y = 16'h200;
			16'h480a: y = 16'h200;
			16'h480b: y = 16'h200;
			16'h480c: y = 16'h200;
			16'h480d: y = 16'h200;
			16'h480e: y = 16'h200;
			16'h480f: y = 16'h200;
			16'h4810: y = 16'h200;
			16'h4811: y = 16'h200;
			16'h4812: y = 16'h200;
			16'h4813: y = 16'h200;
			16'h4814: y = 16'h200;
			16'h4815: y = 16'h200;
			16'h4816: y = 16'h200;
			16'h4817: y = 16'h200;
			16'h4818: y = 16'h200;
			16'h4819: y = 16'h200;
			16'h481a: y = 16'h200;
			16'h481b: y = 16'h200;
			16'h481c: y = 16'h200;
			16'h481d: y = 16'h200;
			16'h481e: y = 16'h200;
			16'h481f: y = 16'h200;
			16'h4820: y = 16'h200;
			16'h4821: y = 16'h200;
			16'h4822: y = 16'h200;
			16'h4823: y = 16'h200;
			16'h4824: y = 16'h200;
			16'h4825: y = 16'h200;
			16'h4826: y = 16'h200;
			16'h4827: y = 16'h200;
			16'h4828: y = 16'h200;
			16'h4829: y = 16'h200;
			16'h482a: y = 16'h200;
			16'h482b: y = 16'h200;
			16'h482c: y = 16'h200;
			16'h482d: y = 16'h200;
			16'h482e: y = 16'h200;
			16'h482f: y = 16'h200;
			16'h4830: y = 16'h200;
			16'h4831: y = 16'h200;
			16'h4832: y = 16'h200;
			16'h4833: y = 16'h200;
			16'h4834: y = 16'h200;
			16'h4835: y = 16'h200;
			16'h4836: y = 16'h200;
			16'h4837: y = 16'h200;
			16'h4838: y = 16'h200;
			16'h4839: y = 16'h200;
			16'h483a: y = 16'h200;
			16'h483b: y = 16'h200;
			16'h483c: y = 16'h200;
			16'h483d: y = 16'h200;
			16'h483e: y = 16'h200;
			16'h483f: y = 16'h200;
			16'h4840: y = 16'h200;
			16'h4841: y = 16'h200;
			16'h4842: y = 16'h200;
			16'h4843: y = 16'h200;
			16'h4844: y = 16'h200;
			16'h4845: y = 16'h200;
			16'h4846: y = 16'h200;
			16'h4847: y = 16'h200;
			16'h4848: y = 16'h200;
			16'h4849: y = 16'h200;
			16'h484a: y = 16'h200;
			16'h484b: y = 16'h200;
			16'h484c: y = 16'h200;
			16'h484d: y = 16'h200;
			16'h484e: y = 16'h200;
			16'h484f: y = 16'h200;
			16'h4850: y = 16'h200;
			16'h4851: y = 16'h200;
			16'h4852: y = 16'h200;
			16'h4853: y = 16'h200;
			16'h4854: y = 16'h200;
			16'h4855: y = 16'h200;
			16'h4856: y = 16'h200;
			16'h4857: y = 16'h200;
			16'h4858: y = 16'h200;
			16'h4859: y = 16'h200;
			16'h485a: y = 16'h200;
			16'h485b: y = 16'h200;
			16'h485c: y = 16'h200;
			16'h485d: y = 16'h200;
			16'h485e: y = 16'h200;
			16'h485f: y = 16'h200;
			16'h4860: y = 16'h200;
			16'h4861: y = 16'h200;
			16'h4862: y = 16'h200;
			16'h4863: y = 16'h200;
			16'h4864: y = 16'h200;
			16'h4865: y = 16'h200;
			16'h4866: y = 16'h200;
			16'h4867: y = 16'h200;
			16'h4868: y = 16'h200;
			16'h4869: y = 16'h200;
			16'h486a: y = 16'h200;
			16'h486b: y = 16'h200;
			16'h486c: y = 16'h200;
			16'h486d: y = 16'h200;
			16'h486e: y = 16'h200;
			16'h486f: y = 16'h200;
			16'h4870: y = 16'h200;
			16'h4871: y = 16'h200;
			16'h4872: y = 16'h200;
			16'h4873: y = 16'h200;
			16'h4874: y = 16'h200;
			16'h4875: y = 16'h200;
			16'h4876: y = 16'h200;
			16'h4877: y = 16'h200;
			16'h4878: y = 16'h200;
			16'h4879: y = 16'h200;
			16'h487a: y = 16'h200;
			16'h487b: y = 16'h200;
			16'h487c: y = 16'h200;
			16'h487d: y = 16'h200;
			16'h487e: y = 16'h200;
			16'h487f: y = 16'h200;
			16'h4880: y = 16'h200;
			16'h4881: y = 16'h200;
			16'h4882: y = 16'h200;
			16'h4883: y = 16'h200;
			16'h4884: y = 16'h200;
			16'h4885: y = 16'h200;
			16'h4886: y = 16'h200;
			16'h4887: y = 16'h200;
			16'h4888: y = 16'h200;
			16'h4889: y = 16'h200;
			16'h488a: y = 16'h200;
			16'h488b: y = 16'h200;
			16'h488c: y = 16'h200;
			16'h488d: y = 16'h200;
			16'h488e: y = 16'h200;
			16'h488f: y = 16'h200;
			16'h4890: y = 16'h200;
			16'h4891: y = 16'h200;
			16'h4892: y = 16'h200;
			16'h4893: y = 16'h200;
			16'h4894: y = 16'h200;
			16'h4895: y = 16'h200;
			16'h4896: y = 16'h200;
			16'h4897: y = 16'h200;
			16'h4898: y = 16'h200;
			16'h4899: y = 16'h200;
			16'h489a: y = 16'h200;
			16'h489b: y = 16'h200;
			16'h489c: y = 16'h200;
			16'h489d: y = 16'h200;
			16'h489e: y = 16'h200;
			16'h489f: y = 16'h200;
			16'h48a0: y = 16'h200;
			16'h48a1: y = 16'h200;
			16'h48a2: y = 16'h200;
			16'h48a3: y = 16'h200;
			16'h48a4: y = 16'h200;
			16'h48a5: y = 16'h200;
			16'h48a6: y = 16'h200;
			16'h48a7: y = 16'h200;
			16'h48a8: y = 16'h200;
			16'h48a9: y = 16'h200;
			16'h48aa: y = 16'h200;
			16'h48ab: y = 16'h200;
			16'h48ac: y = 16'h200;
			16'h48ad: y = 16'h200;
			16'h48ae: y = 16'h200;
			16'h48af: y = 16'h200;
			16'h48b0: y = 16'h200;
			16'h48b1: y = 16'h200;
			16'h48b2: y = 16'h200;
			16'h48b3: y = 16'h200;
			16'h48b4: y = 16'h200;
			16'h48b5: y = 16'h200;
			16'h48b6: y = 16'h200;
			16'h48b7: y = 16'h200;
			16'h48b8: y = 16'h200;
			16'h48b9: y = 16'h200;
			16'h48ba: y = 16'h200;
			16'h48bb: y = 16'h200;
			16'h48bc: y = 16'h200;
			16'h48bd: y = 16'h200;
			16'h48be: y = 16'h200;
			16'h48bf: y = 16'h200;
			16'h48c0: y = 16'h200;
			16'h48c1: y = 16'h200;
			16'h48c2: y = 16'h200;
			16'h48c3: y = 16'h200;
			16'h48c4: y = 16'h200;
			16'h48c5: y = 16'h200;
			16'h48c6: y = 16'h200;
			16'h48c7: y = 16'h200;
			16'h48c8: y = 16'h200;
			16'h48c9: y = 16'h200;
			16'h48ca: y = 16'h200;
			16'h48cb: y = 16'h200;
			16'h48cc: y = 16'h200;
			16'h48cd: y = 16'h200;
			16'h48ce: y = 16'h200;
			16'h48cf: y = 16'h200;
			16'h48d0: y = 16'h200;
			16'h48d1: y = 16'h200;
			16'h48d2: y = 16'h200;
			16'h48d3: y = 16'h200;
			16'h48d4: y = 16'h200;
			16'h48d5: y = 16'h200;
			16'h48d6: y = 16'h200;
			16'h48d7: y = 16'h200;
			16'h48d8: y = 16'h200;
			16'h48d9: y = 16'h200;
			16'h48da: y = 16'h200;
			16'h48db: y = 16'h200;
			16'h48dc: y = 16'h200;
			16'h48dd: y = 16'h200;
			16'h48de: y = 16'h200;
			16'h48df: y = 16'h200;
			16'h48e0: y = 16'h200;
			16'h48e1: y = 16'h200;
			16'h48e2: y = 16'h200;
			16'h48e3: y = 16'h200;
			16'h48e4: y = 16'h200;
			16'h48e5: y = 16'h200;
			16'h48e6: y = 16'h200;
			16'h48e7: y = 16'h200;
			16'h48e8: y = 16'h200;
			16'h48e9: y = 16'h200;
			16'h48ea: y = 16'h200;
			16'h48eb: y = 16'h200;
			16'h48ec: y = 16'h200;
			16'h48ed: y = 16'h200;
			16'h48ee: y = 16'h200;
			16'h48ef: y = 16'h200;
			16'h48f0: y = 16'h200;
			16'h48f1: y = 16'h200;
			16'h48f2: y = 16'h200;
			16'h48f3: y = 16'h200;
			16'h48f4: y = 16'h200;
			16'h48f5: y = 16'h200;
			16'h48f6: y = 16'h200;
			16'h48f7: y = 16'h200;
			16'h48f8: y = 16'h200;
			16'h48f9: y = 16'h200;
			16'h48fa: y = 16'h200;
			16'h48fb: y = 16'h200;
			16'h48fc: y = 16'h200;
			16'h48fd: y = 16'h200;
			16'h48fe: y = 16'h200;
			16'h48ff: y = 16'h200;
			16'h4900: y = 16'h200;
			16'h4901: y = 16'h200;
			16'h4902: y = 16'h200;
			16'h4903: y = 16'h200;
			16'h4904: y = 16'h200;
			16'h4905: y = 16'h200;
			16'h4906: y = 16'h200;
			16'h4907: y = 16'h200;
			16'h4908: y = 16'h200;
			16'h4909: y = 16'h200;
			16'h490a: y = 16'h200;
			16'h490b: y = 16'h200;
			16'h490c: y = 16'h200;
			16'h490d: y = 16'h200;
			16'h490e: y = 16'h200;
			16'h490f: y = 16'h200;
			16'h4910: y = 16'h200;
			16'h4911: y = 16'h200;
			16'h4912: y = 16'h200;
			16'h4913: y = 16'h200;
			16'h4914: y = 16'h200;
			16'h4915: y = 16'h200;
			16'h4916: y = 16'h200;
			16'h4917: y = 16'h200;
			16'h4918: y = 16'h200;
			16'h4919: y = 16'h200;
			16'h491a: y = 16'h200;
			16'h491b: y = 16'h200;
			16'h491c: y = 16'h200;
			16'h491d: y = 16'h200;
			16'h491e: y = 16'h200;
			16'h491f: y = 16'h200;
			16'h4920: y = 16'h200;
			16'h4921: y = 16'h200;
			16'h4922: y = 16'h200;
			16'h4923: y = 16'h200;
			16'h4924: y = 16'h200;
			16'h4925: y = 16'h200;
			16'h4926: y = 16'h200;
			16'h4927: y = 16'h200;
			16'h4928: y = 16'h200;
			16'h4929: y = 16'h200;
			16'h492a: y = 16'h200;
			16'h492b: y = 16'h200;
			16'h492c: y = 16'h200;
			16'h492d: y = 16'h200;
			16'h492e: y = 16'h200;
			16'h492f: y = 16'h200;
			16'h4930: y = 16'h200;
			16'h4931: y = 16'h200;
			16'h4932: y = 16'h200;
			16'h4933: y = 16'h200;
			16'h4934: y = 16'h200;
			16'h4935: y = 16'h200;
			16'h4936: y = 16'h200;
			16'h4937: y = 16'h200;
			16'h4938: y = 16'h200;
			16'h4939: y = 16'h200;
			16'h493a: y = 16'h200;
			16'h493b: y = 16'h200;
			16'h493c: y = 16'h200;
			16'h493d: y = 16'h200;
			16'h493e: y = 16'h200;
			16'h493f: y = 16'h200;
			16'h4940: y = 16'h200;
			16'h4941: y = 16'h200;
			16'h4942: y = 16'h200;
			16'h4943: y = 16'h200;
			16'h4944: y = 16'h200;
			16'h4945: y = 16'h200;
			16'h4946: y = 16'h200;
			16'h4947: y = 16'h200;
			16'h4948: y = 16'h200;
			16'h4949: y = 16'h200;
			16'h494a: y = 16'h200;
			16'h494b: y = 16'h200;
			16'h494c: y = 16'h200;
			16'h494d: y = 16'h200;
			16'h494e: y = 16'h200;
			16'h494f: y = 16'h200;
			16'h4950: y = 16'h200;
			16'h4951: y = 16'h200;
			16'h4952: y = 16'h200;
			16'h4953: y = 16'h200;
			16'h4954: y = 16'h200;
			16'h4955: y = 16'h200;
			16'h4956: y = 16'h200;
			16'h4957: y = 16'h200;
			16'h4958: y = 16'h200;
			16'h4959: y = 16'h200;
			16'h495a: y = 16'h200;
			16'h495b: y = 16'h200;
			16'h495c: y = 16'h200;
			16'h495d: y = 16'h200;
			16'h495e: y = 16'h200;
			16'h495f: y = 16'h200;
			16'h4960: y = 16'h200;
			16'h4961: y = 16'h200;
			16'h4962: y = 16'h200;
			16'h4963: y = 16'h200;
			16'h4964: y = 16'h200;
			16'h4965: y = 16'h200;
			16'h4966: y = 16'h200;
			16'h4967: y = 16'h200;
			16'h4968: y = 16'h200;
			16'h4969: y = 16'h200;
			16'h496a: y = 16'h200;
			16'h496b: y = 16'h200;
			16'h496c: y = 16'h200;
			16'h496d: y = 16'h200;
			16'h496e: y = 16'h200;
			16'h496f: y = 16'h200;
			16'h4970: y = 16'h200;
			16'h4971: y = 16'h200;
			16'h4972: y = 16'h200;
			16'h4973: y = 16'h200;
			16'h4974: y = 16'h200;
			16'h4975: y = 16'h200;
			16'h4976: y = 16'h200;
			16'h4977: y = 16'h200;
			16'h4978: y = 16'h200;
			16'h4979: y = 16'h200;
			16'h497a: y = 16'h200;
			16'h497b: y = 16'h200;
			16'h497c: y = 16'h200;
			16'h497d: y = 16'h200;
			16'h497e: y = 16'h200;
			16'h497f: y = 16'h200;
			16'h4980: y = 16'h200;
			16'h4981: y = 16'h200;
			16'h4982: y = 16'h200;
			16'h4983: y = 16'h200;
			16'h4984: y = 16'h200;
			16'h4985: y = 16'h200;
			16'h4986: y = 16'h200;
			16'h4987: y = 16'h200;
			16'h4988: y = 16'h200;
			16'h4989: y = 16'h200;
			16'h498a: y = 16'h200;
			16'h498b: y = 16'h200;
			16'h498c: y = 16'h200;
			16'h498d: y = 16'h200;
			16'h498e: y = 16'h200;
			16'h498f: y = 16'h200;
			16'h4990: y = 16'h200;
			16'h4991: y = 16'h200;
			16'h4992: y = 16'h200;
			16'h4993: y = 16'h200;
			16'h4994: y = 16'h200;
			16'h4995: y = 16'h200;
			16'h4996: y = 16'h200;
			16'h4997: y = 16'h200;
			16'h4998: y = 16'h200;
			16'h4999: y = 16'h200;
			16'h499a: y = 16'h200;
			16'h499b: y = 16'h200;
			16'h499c: y = 16'h200;
			16'h499d: y = 16'h200;
			16'h499e: y = 16'h200;
			16'h499f: y = 16'h200;
			16'h49a0: y = 16'h200;
			16'h49a1: y = 16'h200;
			16'h49a2: y = 16'h200;
			16'h49a3: y = 16'h200;
			16'h49a4: y = 16'h200;
			16'h49a5: y = 16'h200;
			16'h49a6: y = 16'h200;
			16'h49a7: y = 16'h200;
			16'h49a8: y = 16'h200;
			16'h49a9: y = 16'h200;
			16'h49aa: y = 16'h200;
			16'h49ab: y = 16'h200;
			16'h49ac: y = 16'h200;
			16'h49ad: y = 16'h200;
			16'h49ae: y = 16'h200;
			16'h49af: y = 16'h200;
			16'h49b0: y = 16'h200;
			16'h49b1: y = 16'h200;
			16'h49b2: y = 16'h200;
			16'h49b3: y = 16'h200;
			16'h49b4: y = 16'h200;
			16'h49b5: y = 16'h200;
			16'h49b6: y = 16'h200;
			16'h49b7: y = 16'h200;
			16'h49b8: y = 16'h200;
			16'h49b9: y = 16'h200;
			16'h49ba: y = 16'h200;
			16'h49bb: y = 16'h200;
			16'h49bc: y = 16'h200;
			16'h49bd: y = 16'h200;
			16'h49be: y = 16'h200;
			16'h49bf: y = 16'h200;
			16'h49c0: y = 16'h200;
			16'h49c1: y = 16'h200;
			16'h49c2: y = 16'h200;
			16'h49c3: y = 16'h200;
			16'h49c4: y = 16'h200;
			16'h49c5: y = 16'h200;
			16'h49c6: y = 16'h200;
			16'h49c7: y = 16'h200;
			16'h49c8: y = 16'h200;
			16'h49c9: y = 16'h200;
			16'h49ca: y = 16'h200;
			16'h49cb: y = 16'h200;
			16'h49cc: y = 16'h200;
			16'h49cd: y = 16'h200;
			16'h49ce: y = 16'h200;
			16'h49cf: y = 16'h200;
			16'h49d0: y = 16'h200;
			16'h49d1: y = 16'h200;
			16'h49d2: y = 16'h200;
			16'h49d3: y = 16'h200;
			16'h49d4: y = 16'h200;
			16'h49d5: y = 16'h200;
			16'h49d6: y = 16'h200;
			16'h49d7: y = 16'h200;
			16'h49d8: y = 16'h200;
			16'h49d9: y = 16'h200;
			16'h49da: y = 16'h200;
			16'h49db: y = 16'h200;
			16'h49dc: y = 16'h200;
			16'h49dd: y = 16'h200;
			16'h49de: y = 16'h200;
			16'h49df: y = 16'h200;
			16'h49e0: y = 16'h200;
			16'h49e1: y = 16'h200;
			16'h49e2: y = 16'h200;
			16'h49e3: y = 16'h200;
			16'h49e4: y = 16'h200;
			16'h49e5: y = 16'h200;
			16'h49e6: y = 16'h200;
			16'h49e7: y = 16'h200;
			16'h49e8: y = 16'h200;
			16'h49e9: y = 16'h200;
			16'h49ea: y = 16'h200;
			16'h49eb: y = 16'h200;
			16'h49ec: y = 16'h200;
			16'h49ed: y = 16'h200;
			16'h49ee: y = 16'h200;
			16'h49ef: y = 16'h200;
			16'h49f0: y = 16'h200;
			16'h49f1: y = 16'h200;
			16'h49f2: y = 16'h200;
			16'h49f3: y = 16'h200;
			16'h49f4: y = 16'h200;
			16'h49f5: y = 16'h200;
			16'h49f6: y = 16'h200;
			16'h49f7: y = 16'h200;
			16'h49f8: y = 16'h200;
			16'h49f9: y = 16'h200;
			16'h49fa: y = 16'h200;
			16'h49fb: y = 16'h200;
			16'h49fc: y = 16'h200;
			16'h49fd: y = 16'h200;
			16'h49fe: y = 16'h200;
			16'h49ff: y = 16'h200;
			16'h4a00: y = 16'h200;
			16'h4a01: y = 16'h200;
			16'h4a02: y = 16'h200;
			16'h4a03: y = 16'h200;
			16'h4a04: y = 16'h200;
			16'h4a05: y = 16'h200;
			16'h4a06: y = 16'h200;
			16'h4a07: y = 16'h200;
			16'h4a08: y = 16'h200;
			16'h4a09: y = 16'h200;
			16'h4a0a: y = 16'h200;
			16'h4a0b: y = 16'h200;
			16'h4a0c: y = 16'h200;
			16'h4a0d: y = 16'h200;
			16'h4a0e: y = 16'h200;
			16'h4a0f: y = 16'h200;
			16'h4a10: y = 16'h200;
			16'h4a11: y = 16'h200;
			16'h4a12: y = 16'h200;
			16'h4a13: y = 16'h200;
			16'h4a14: y = 16'h200;
			16'h4a15: y = 16'h200;
			16'h4a16: y = 16'h200;
			16'h4a17: y = 16'h200;
			16'h4a18: y = 16'h200;
			16'h4a19: y = 16'h200;
			16'h4a1a: y = 16'h200;
			16'h4a1b: y = 16'h200;
			16'h4a1c: y = 16'h200;
			16'h4a1d: y = 16'h200;
			16'h4a1e: y = 16'h200;
			16'h4a1f: y = 16'h200;
			16'h4a20: y = 16'h200;
			16'h4a21: y = 16'h200;
			16'h4a22: y = 16'h200;
			16'h4a23: y = 16'h200;
			16'h4a24: y = 16'h200;
			16'h4a25: y = 16'h200;
			16'h4a26: y = 16'h200;
			16'h4a27: y = 16'h200;
			16'h4a28: y = 16'h200;
			16'h4a29: y = 16'h200;
			16'h4a2a: y = 16'h200;
			16'h4a2b: y = 16'h200;
			16'h4a2c: y = 16'h200;
			16'h4a2d: y = 16'h200;
			16'h4a2e: y = 16'h200;
			16'h4a2f: y = 16'h200;
			16'h4a30: y = 16'h200;
			16'h4a31: y = 16'h200;
			16'h4a32: y = 16'h200;
			16'h4a33: y = 16'h200;
			16'h4a34: y = 16'h200;
			16'h4a35: y = 16'h200;
			16'h4a36: y = 16'h200;
			16'h4a37: y = 16'h200;
			16'h4a38: y = 16'h200;
			16'h4a39: y = 16'h200;
			16'h4a3a: y = 16'h200;
			16'h4a3b: y = 16'h200;
			16'h4a3c: y = 16'h200;
			16'h4a3d: y = 16'h200;
			16'h4a3e: y = 16'h200;
			16'h4a3f: y = 16'h200;
			16'h4a40: y = 16'h200;
			16'h4a41: y = 16'h200;
			16'h4a42: y = 16'h200;
			16'h4a43: y = 16'h200;
			16'h4a44: y = 16'h200;
			16'h4a45: y = 16'h200;
			16'h4a46: y = 16'h200;
			16'h4a47: y = 16'h200;
			16'h4a48: y = 16'h200;
			16'h4a49: y = 16'h200;
			16'h4a4a: y = 16'h200;
			16'h4a4b: y = 16'h200;
			16'h4a4c: y = 16'h200;
			16'h4a4d: y = 16'h200;
			16'h4a4e: y = 16'h200;
			16'h4a4f: y = 16'h200;
			16'h4a50: y = 16'h200;
			16'h4a51: y = 16'h200;
			16'h4a52: y = 16'h200;
			16'h4a53: y = 16'h200;
			16'h4a54: y = 16'h200;
			16'h4a55: y = 16'h200;
			16'h4a56: y = 16'h200;
			16'h4a57: y = 16'h200;
			16'h4a58: y = 16'h200;
			16'h4a59: y = 16'h200;
			16'h4a5a: y = 16'h200;
			16'h4a5b: y = 16'h200;
			16'h4a5c: y = 16'h200;
			16'h4a5d: y = 16'h200;
			16'h4a5e: y = 16'h200;
			16'h4a5f: y = 16'h200;
			16'h4a60: y = 16'h200;
			16'h4a61: y = 16'h200;
			16'h4a62: y = 16'h200;
			16'h4a63: y = 16'h200;
			16'h4a64: y = 16'h200;
			16'h4a65: y = 16'h200;
			16'h4a66: y = 16'h200;
			16'h4a67: y = 16'h200;
			16'h4a68: y = 16'h200;
			16'h4a69: y = 16'h200;
			16'h4a6a: y = 16'h200;
			16'h4a6b: y = 16'h200;
			16'h4a6c: y = 16'h200;
			16'h4a6d: y = 16'h200;
			16'h4a6e: y = 16'h200;
			16'h4a6f: y = 16'h200;
			16'h4a70: y = 16'h200;
			16'h4a71: y = 16'h200;
			16'h4a72: y = 16'h200;
			16'h4a73: y = 16'h200;
			16'h4a74: y = 16'h200;
			16'h4a75: y = 16'h200;
			16'h4a76: y = 16'h200;
			16'h4a77: y = 16'h200;
			16'h4a78: y = 16'h200;
			16'h4a79: y = 16'h200;
			16'h4a7a: y = 16'h200;
			16'h4a7b: y = 16'h200;
			16'h4a7c: y = 16'h200;
			16'h4a7d: y = 16'h200;
			16'h4a7e: y = 16'h200;
			16'h4a7f: y = 16'h200;
			16'h4a80: y = 16'h200;
			16'h4a81: y = 16'h200;
			16'h4a82: y = 16'h200;
			16'h4a83: y = 16'h200;
			16'h4a84: y = 16'h200;
			16'h4a85: y = 16'h200;
			16'h4a86: y = 16'h200;
			16'h4a87: y = 16'h200;
			16'h4a88: y = 16'h200;
			16'h4a89: y = 16'h200;
			16'h4a8a: y = 16'h200;
			16'h4a8b: y = 16'h200;
			16'h4a8c: y = 16'h200;
			16'h4a8d: y = 16'h200;
			16'h4a8e: y = 16'h200;
			16'h4a8f: y = 16'h200;
			16'h4a90: y = 16'h200;
			16'h4a91: y = 16'h200;
			16'h4a92: y = 16'h200;
			16'h4a93: y = 16'h200;
			16'h4a94: y = 16'h200;
			16'h4a95: y = 16'h200;
			16'h4a96: y = 16'h200;
			16'h4a97: y = 16'h200;
			16'h4a98: y = 16'h200;
			16'h4a99: y = 16'h200;
			16'h4a9a: y = 16'h200;
			16'h4a9b: y = 16'h200;
			16'h4a9c: y = 16'h200;
			16'h4a9d: y = 16'h200;
			16'h4a9e: y = 16'h200;
			16'h4a9f: y = 16'h200;
			16'h4aa0: y = 16'h200;
			16'h4aa1: y = 16'h200;
			16'h4aa2: y = 16'h200;
			16'h4aa3: y = 16'h200;
			16'h4aa4: y = 16'h200;
			16'h4aa5: y = 16'h200;
			16'h4aa6: y = 16'h200;
			16'h4aa7: y = 16'h200;
			16'h4aa8: y = 16'h200;
			16'h4aa9: y = 16'h200;
			16'h4aaa: y = 16'h200;
			16'h4aab: y = 16'h200;
			16'h4aac: y = 16'h200;
			16'h4aad: y = 16'h200;
			16'h4aae: y = 16'h200;
			16'h4aaf: y = 16'h200;
			16'h4ab0: y = 16'h200;
			16'h4ab1: y = 16'h200;
			16'h4ab2: y = 16'h200;
			16'h4ab3: y = 16'h200;
			16'h4ab4: y = 16'h200;
			16'h4ab5: y = 16'h200;
			16'h4ab6: y = 16'h200;
			16'h4ab7: y = 16'h200;
			16'h4ab8: y = 16'h200;
			16'h4ab9: y = 16'h200;
			16'h4aba: y = 16'h200;
			16'h4abb: y = 16'h200;
			16'h4abc: y = 16'h200;
			16'h4abd: y = 16'h200;
			16'h4abe: y = 16'h200;
			16'h4abf: y = 16'h200;
			16'h4ac0: y = 16'h200;
			16'h4ac1: y = 16'h200;
			16'h4ac2: y = 16'h200;
			16'h4ac3: y = 16'h200;
			16'h4ac4: y = 16'h200;
			16'h4ac5: y = 16'h200;
			16'h4ac6: y = 16'h200;
			16'h4ac7: y = 16'h200;
			16'h4ac8: y = 16'h200;
			16'h4ac9: y = 16'h200;
			16'h4aca: y = 16'h200;
			16'h4acb: y = 16'h200;
			16'h4acc: y = 16'h200;
			16'h4acd: y = 16'h200;
			16'h4ace: y = 16'h200;
			16'h4acf: y = 16'h200;
			16'h4ad0: y = 16'h200;
			16'h4ad1: y = 16'h200;
			16'h4ad2: y = 16'h200;
			16'h4ad3: y = 16'h200;
			16'h4ad4: y = 16'h200;
			16'h4ad5: y = 16'h200;
			16'h4ad6: y = 16'h200;
			16'h4ad7: y = 16'h200;
			16'h4ad8: y = 16'h200;
			16'h4ad9: y = 16'h200;
			16'h4ada: y = 16'h200;
			16'h4adb: y = 16'h200;
			16'h4adc: y = 16'h200;
			16'h4add: y = 16'h200;
			16'h4ade: y = 16'h200;
			16'h4adf: y = 16'h200;
			16'h4ae0: y = 16'h200;
			16'h4ae1: y = 16'h200;
			16'h4ae2: y = 16'h200;
			16'h4ae3: y = 16'h200;
			16'h4ae4: y = 16'h200;
			16'h4ae5: y = 16'h200;
			16'h4ae6: y = 16'h200;
			16'h4ae7: y = 16'h200;
			16'h4ae8: y = 16'h200;
			16'h4ae9: y = 16'h200;
			16'h4aea: y = 16'h200;
			16'h4aeb: y = 16'h200;
			16'h4aec: y = 16'h200;
			16'h4aed: y = 16'h200;
			16'h4aee: y = 16'h200;
			16'h4aef: y = 16'h200;
			16'h4af0: y = 16'h200;
			16'h4af1: y = 16'h200;
			16'h4af2: y = 16'h200;
			16'h4af3: y = 16'h200;
			16'h4af4: y = 16'h200;
			16'h4af5: y = 16'h200;
			16'h4af6: y = 16'h200;
			16'h4af7: y = 16'h200;
			16'h4af8: y = 16'h200;
			16'h4af9: y = 16'h200;
			16'h4afa: y = 16'h200;
			16'h4afb: y = 16'h200;
			16'h4afc: y = 16'h200;
			16'h4afd: y = 16'h200;
			16'h4afe: y = 16'h200;
			16'h4aff: y = 16'h200;
			16'h4b00: y = 16'h200;
			16'h4b01: y = 16'h200;
			16'h4b02: y = 16'h200;
			16'h4b03: y = 16'h200;
			16'h4b04: y = 16'h200;
			16'h4b05: y = 16'h200;
			16'h4b06: y = 16'h200;
			16'h4b07: y = 16'h200;
			16'h4b08: y = 16'h200;
			16'h4b09: y = 16'h200;
			16'h4b0a: y = 16'h200;
			16'h4b0b: y = 16'h200;
			16'h4b0c: y = 16'h200;
			16'h4b0d: y = 16'h200;
			16'h4b0e: y = 16'h200;
			16'h4b0f: y = 16'h200;
			16'h4b10: y = 16'h200;
			16'h4b11: y = 16'h200;
			16'h4b12: y = 16'h200;
			16'h4b13: y = 16'h200;
			16'h4b14: y = 16'h200;
			16'h4b15: y = 16'h200;
			16'h4b16: y = 16'h200;
			16'h4b17: y = 16'h200;
			16'h4b18: y = 16'h200;
			16'h4b19: y = 16'h200;
			16'h4b1a: y = 16'h200;
			16'h4b1b: y = 16'h200;
			16'h4b1c: y = 16'h200;
			16'h4b1d: y = 16'h200;
			16'h4b1e: y = 16'h200;
			16'h4b1f: y = 16'h200;
			16'h4b20: y = 16'h200;
			16'h4b21: y = 16'h200;
			16'h4b22: y = 16'h200;
			16'h4b23: y = 16'h200;
			16'h4b24: y = 16'h200;
			16'h4b25: y = 16'h200;
			16'h4b26: y = 16'h200;
			16'h4b27: y = 16'h200;
			16'h4b28: y = 16'h200;
			16'h4b29: y = 16'h200;
			16'h4b2a: y = 16'h200;
			16'h4b2b: y = 16'h200;
			16'h4b2c: y = 16'h200;
			16'h4b2d: y = 16'h200;
			16'h4b2e: y = 16'h200;
			16'h4b2f: y = 16'h200;
			16'h4b30: y = 16'h200;
			16'h4b31: y = 16'h200;
			16'h4b32: y = 16'h200;
			16'h4b33: y = 16'h200;
			16'h4b34: y = 16'h200;
			16'h4b35: y = 16'h200;
			16'h4b36: y = 16'h200;
			16'h4b37: y = 16'h200;
			16'h4b38: y = 16'h200;
			16'h4b39: y = 16'h200;
			16'h4b3a: y = 16'h200;
			16'h4b3b: y = 16'h200;
			16'h4b3c: y = 16'h200;
			16'h4b3d: y = 16'h200;
			16'h4b3e: y = 16'h200;
			16'h4b3f: y = 16'h200;
			16'h4b40: y = 16'h200;
			16'h4b41: y = 16'h200;
			16'h4b42: y = 16'h200;
			16'h4b43: y = 16'h200;
			16'h4b44: y = 16'h200;
			16'h4b45: y = 16'h200;
			16'h4b46: y = 16'h200;
			16'h4b47: y = 16'h200;
			16'h4b48: y = 16'h200;
			16'h4b49: y = 16'h200;
			16'h4b4a: y = 16'h200;
			16'h4b4b: y = 16'h200;
			16'h4b4c: y = 16'h200;
			16'h4b4d: y = 16'h200;
			16'h4b4e: y = 16'h200;
			16'h4b4f: y = 16'h200;
			16'h4b50: y = 16'h200;
			16'h4b51: y = 16'h200;
			16'h4b52: y = 16'h200;
			16'h4b53: y = 16'h200;
			16'h4b54: y = 16'h200;
			16'h4b55: y = 16'h200;
			16'h4b56: y = 16'h200;
			16'h4b57: y = 16'h200;
			16'h4b58: y = 16'h200;
			16'h4b59: y = 16'h200;
			16'h4b5a: y = 16'h200;
			16'h4b5b: y = 16'h200;
			16'h4b5c: y = 16'h200;
			16'h4b5d: y = 16'h200;
			16'h4b5e: y = 16'h200;
			16'h4b5f: y = 16'h200;
			16'h4b60: y = 16'h200;
			16'h4b61: y = 16'h200;
			16'h4b62: y = 16'h200;
			16'h4b63: y = 16'h200;
			16'h4b64: y = 16'h200;
			16'h4b65: y = 16'h200;
			16'h4b66: y = 16'h200;
			16'h4b67: y = 16'h200;
			16'h4b68: y = 16'h200;
			16'h4b69: y = 16'h200;
			16'h4b6a: y = 16'h200;
			16'h4b6b: y = 16'h200;
			16'h4b6c: y = 16'h200;
			16'h4b6d: y = 16'h200;
			16'h4b6e: y = 16'h200;
			16'h4b6f: y = 16'h200;
			16'h4b70: y = 16'h200;
			16'h4b71: y = 16'h200;
			16'h4b72: y = 16'h200;
			16'h4b73: y = 16'h200;
			16'h4b74: y = 16'h200;
			16'h4b75: y = 16'h200;
			16'h4b76: y = 16'h200;
			16'h4b77: y = 16'h200;
			16'h4b78: y = 16'h200;
			16'h4b79: y = 16'h200;
			16'h4b7a: y = 16'h200;
			16'h4b7b: y = 16'h200;
			16'h4b7c: y = 16'h200;
			16'h4b7d: y = 16'h200;
			16'h4b7e: y = 16'h200;
			16'h4b7f: y = 16'h200;
			16'h4b80: y = 16'h200;
			16'h4b81: y = 16'h200;
			16'h4b82: y = 16'h200;
			16'h4b83: y = 16'h200;
			16'h4b84: y = 16'h200;
			16'h4b85: y = 16'h200;
			16'h4b86: y = 16'h200;
			16'h4b87: y = 16'h200;
			16'h4b88: y = 16'h200;
			16'h4b89: y = 16'h200;
			16'h4b8a: y = 16'h200;
			16'h4b8b: y = 16'h200;
			16'h4b8c: y = 16'h200;
			16'h4b8d: y = 16'h200;
			16'h4b8e: y = 16'h200;
			16'h4b8f: y = 16'h200;
			16'h4b90: y = 16'h200;
			16'h4b91: y = 16'h200;
			16'h4b92: y = 16'h200;
			16'h4b93: y = 16'h200;
			16'h4b94: y = 16'h200;
			16'h4b95: y = 16'h200;
			16'h4b96: y = 16'h200;
			16'h4b97: y = 16'h200;
			16'h4b98: y = 16'h200;
			16'h4b99: y = 16'h200;
			16'h4b9a: y = 16'h200;
			16'h4b9b: y = 16'h200;
			16'h4b9c: y = 16'h200;
			16'h4b9d: y = 16'h200;
			16'h4b9e: y = 16'h200;
			16'h4b9f: y = 16'h200;
			16'h4ba0: y = 16'h200;
			16'h4ba1: y = 16'h200;
			16'h4ba2: y = 16'h200;
			16'h4ba3: y = 16'h200;
			16'h4ba4: y = 16'h200;
			16'h4ba5: y = 16'h200;
			16'h4ba6: y = 16'h200;
			16'h4ba7: y = 16'h200;
			16'h4ba8: y = 16'h200;
			16'h4ba9: y = 16'h200;
			16'h4baa: y = 16'h200;
			16'h4bab: y = 16'h200;
			16'h4bac: y = 16'h200;
			16'h4bad: y = 16'h200;
			16'h4bae: y = 16'h200;
			16'h4baf: y = 16'h200;
			16'h4bb0: y = 16'h200;
			16'h4bb1: y = 16'h200;
			16'h4bb2: y = 16'h200;
			16'h4bb3: y = 16'h200;
			16'h4bb4: y = 16'h200;
			16'h4bb5: y = 16'h200;
			16'h4bb6: y = 16'h200;
			16'h4bb7: y = 16'h200;
			16'h4bb8: y = 16'h200;
			16'h4bb9: y = 16'h200;
			16'h4bba: y = 16'h200;
			16'h4bbb: y = 16'h200;
			16'h4bbc: y = 16'h200;
			16'h4bbd: y = 16'h200;
			16'h4bbe: y = 16'h200;
			16'h4bbf: y = 16'h200;
			16'h4bc0: y = 16'h200;
			16'h4bc1: y = 16'h200;
			16'h4bc2: y = 16'h200;
			16'h4bc3: y = 16'h200;
			16'h4bc4: y = 16'h200;
			16'h4bc5: y = 16'h200;
			16'h4bc6: y = 16'h200;
			16'h4bc7: y = 16'h200;
			16'h4bc8: y = 16'h200;
			16'h4bc9: y = 16'h200;
			16'h4bca: y = 16'h200;
			16'h4bcb: y = 16'h200;
			16'h4bcc: y = 16'h200;
			16'h4bcd: y = 16'h200;
			16'h4bce: y = 16'h200;
			16'h4bcf: y = 16'h200;
			16'h4bd0: y = 16'h200;
			16'h4bd1: y = 16'h200;
			16'h4bd2: y = 16'h200;
			16'h4bd3: y = 16'h200;
			16'h4bd4: y = 16'h200;
			16'h4bd5: y = 16'h200;
			16'h4bd6: y = 16'h200;
			16'h4bd7: y = 16'h200;
			16'h4bd8: y = 16'h200;
			16'h4bd9: y = 16'h200;
			16'h4bda: y = 16'h200;
			16'h4bdb: y = 16'h200;
			16'h4bdc: y = 16'h200;
			16'h4bdd: y = 16'h200;
			16'h4bde: y = 16'h200;
			16'h4bdf: y = 16'h200;
			16'h4be0: y = 16'h200;
			16'h4be1: y = 16'h200;
			16'h4be2: y = 16'h200;
			16'h4be3: y = 16'h200;
			16'h4be4: y = 16'h200;
			16'h4be5: y = 16'h200;
			16'h4be6: y = 16'h200;
			16'h4be7: y = 16'h200;
			16'h4be8: y = 16'h200;
			16'h4be9: y = 16'h200;
			16'h4bea: y = 16'h200;
			16'h4beb: y = 16'h200;
			16'h4bec: y = 16'h200;
			16'h4bed: y = 16'h200;
			16'h4bee: y = 16'h200;
			16'h4bef: y = 16'h200;
			16'h4bf0: y = 16'h200;
			16'h4bf1: y = 16'h200;
			16'h4bf2: y = 16'h200;
			16'h4bf3: y = 16'h200;
			16'h4bf4: y = 16'h200;
			16'h4bf5: y = 16'h200;
			16'h4bf6: y = 16'h200;
			16'h4bf7: y = 16'h200;
			16'h4bf8: y = 16'h200;
			16'h4bf9: y = 16'h200;
			16'h4bfa: y = 16'h200;
			16'h4bfb: y = 16'h200;
			16'h4bfc: y = 16'h200;
			16'h4bfd: y = 16'h200;
			16'h4bfe: y = 16'h200;
			16'h4bff: y = 16'h200;
			16'h4c00: y = 16'h200;
			16'h4c01: y = 16'h200;
			16'h4c02: y = 16'h200;
			16'h4c03: y = 16'h200;
			16'h4c04: y = 16'h200;
			16'h4c05: y = 16'h200;
			16'h4c06: y = 16'h200;
			16'h4c07: y = 16'h200;
			16'h4c08: y = 16'h200;
			16'h4c09: y = 16'h200;
			16'h4c0a: y = 16'h200;
			16'h4c0b: y = 16'h200;
			16'h4c0c: y = 16'h200;
			16'h4c0d: y = 16'h200;
			16'h4c0e: y = 16'h200;
			16'h4c0f: y = 16'h200;
			16'h4c10: y = 16'h200;
			16'h4c11: y = 16'h200;
			16'h4c12: y = 16'h200;
			16'h4c13: y = 16'h200;
			16'h4c14: y = 16'h200;
			16'h4c15: y = 16'h200;
			16'h4c16: y = 16'h200;
			16'h4c17: y = 16'h200;
			16'h4c18: y = 16'h200;
			16'h4c19: y = 16'h200;
			16'h4c1a: y = 16'h200;
			16'h4c1b: y = 16'h200;
			16'h4c1c: y = 16'h200;
			16'h4c1d: y = 16'h200;
			16'h4c1e: y = 16'h200;
			16'h4c1f: y = 16'h200;
			16'h4c20: y = 16'h200;
			16'h4c21: y = 16'h200;
			16'h4c22: y = 16'h200;
			16'h4c23: y = 16'h200;
			16'h4c24: y = 16'h200;
			16'h4c25: y = 16'h200;
			16'h4c26: y = 16'h200;
			16'h4c27: y = 16'h200;
			16'h4c28: y = 16'h200;
			16'h4c29: y = 16'h200;
			16'h4c2a: y = 16'h200;
			16'h4c2b: y = 16'h200;
			16'h4c2c: y = 16'h200;
			16'h4c2d: y = 16'h200;
			16'h4c2e: y = 16'h200;
			16'h4c2f: y = 16'h200;
			16'h4c30: y = 16'h200;
			16'h4c31: y = 16'h200;
			16'h4c32: y = 16'h200;
			16'h4c33: y = 16'h200;
			16'h4c34: y = 16'h200;
			16'h4c35: y = 16'h200;
			16'h4c36: y = 16'h200;
			16'h4c37: y = 16'h200;
			16'h4c38: y = 16'h200;
			16'h4c39: y = 16'h200;
			16'h4c3a: y = 16'h200;
			16'h4c3b: y = 16'h200;
			16'h4c3c: y = 16'h200;
			16'h4c3d: y = 16'h200;
			16'h4c3e: y = 16'h200;
			16'h4c3f: y = 16'h200;
			16'h4c40: y = 16'h200;
			16'h4c41: y = 16'h200;
			16'h4c42: y = 16'h200;
			16'h4c43: y = 16'h200;
			16'h4c44: y = 16'h200;
			16'h4c45: y = 16'h200;
			16'h4c46: y = 16'h200;
			16'h4c47: y = 16'h200;
			16'h4c48: y = 16'h200;
			16'h4c49: y = 16'h200;
			16'h4c4a: y = 16'h200;
			16'h4c4b: y = 16'h200;
			16'h4c4c: y = 16'h200;
			16'h4c4d: y = 16'h200;
			16'h4c4e: y = 16'h200;
			16'h4c4f: y = 16'h200;
			16'h4c50: y = 16'h200;
			16'h4c51: y = 16'h200;
			16'h4c52: y = 16'h200;
			16'h4c53: y = 16'h200;
			16'h4c54: y = 16'h200;
			16'h4c55: y = 16'h200;
			16'h4c56: y = 16'h200;
			16'h4c57: y = 16'h200;
			16'h4c58: y = 16'h200;
			16'h4c59: y = 16'h200;
			16'h4c5a: y = 16'h200;
			16'h4c5b: y = 16'h200;
			16'h4c5c: y = 16'h200;
			16'h4c5d: y = 16'h200;
			16'h4c5e: y = 16'h200;
			16'h4c5f: y = 16'h200;
			16'h4c60: y = 16'h200;
			16'h4c61: y = 16'h200;
			16'h4c62: y = 16'h200;
			16'h4c63: y = 16'h200;
			16'h4c64: y = 16'h200;
			16'h4c65: y = 16'h200;
			16'h4c66: y = 16'h200;
			16'h4c67: y = 16'h200;
			16'h4c68: y = 16'h200;
			16'h4c69: y = 16'h200;
			16'h4c6a: y = 16'h200;
			16'h4c6b: y = 16'h200;
			16'h4c6c: y = 16'h200;
			16'h4c6d: y = 16'h200;
			16'h4c6e: y = 16'h200;
			16'h4c6f: y = 16'h200;
			16'h4c70: y = 16'h200;
			16'h4c71: y = 16'h200;
			16'h4c72: y = 16'h200;
			16'h4c73: y = 16'h200;
			16'h4c74: y = 16'h200;
			16'h4c75: y = 16'h200;
			16'h4c76: y = 16'h200;
			16'h4c77: y = 16'h200;
			16'h4c78: y = 16'h200;
			16'h4c79: y = 16'h200;
			16'h4c7a: y = 16'h200;
			16'h4c7b: y = 16'h200;
			16'h4c7c: y = 16'h200;
			16'h4c7d: y = 16'h200;
			16'h4c7e: y = 16'h200;
			16'h4c7f: y = 16'h200;
			16'h4c80: y = 16'h200;
			16'h4c81: y = 16'h200;
			16'h4c82: y = 16'h200;
			16'h4c83: y = 16'h200;
			16'h4c84: y = 16'h200;
			16'h4c85: y = 16'h200;
			16'h4c86: y = 16'h200;
			16'h4c87: y = 16'h200;
			16'h4c88: y = 16'h200;
			16'h4c89: y = 16'h200;
			16'h4c8a: y = 16'h200;
			16'h4c8b: y = 16'h200;
			16'h4c8c: y = 16'h200;
			16'h4c8d: y = 16'h200;
			16'h4c8e: y = 16'h200;
			16'h4c8f: y = 16'h200;
			16'h4c90: y = 16'h200;
			16'h4c91: y = 16'h200;
			16'h4c92: y = 16'h200;
			16'h4c93: y = 16'h200;
			16'h4c94: y = 16'h200;
			16'h4c95: y = 16'h200;
			16'h4c96: y = 16'h200;
			16'h4c97: y = 16'h200;
			16'h4c98: y = 16'h200;
			16'h4c99: y = 16'h200;
			16'h4c9a: y = 16'h200;
			16'h4c9b: y = 16'h200;
			16'h4c9c: y = 16'h200;
			16'h4c9d: y = 16'h200;
			16'h4c9e: y = 16'h200;
			16'h4c9f: y = 16'h200;
			16'h4ca0: y = 16'h200;
			16'h4ca1: y = 16'h200;
			16'h4ca2: y = 16'h200;
			16'h4ca3: y = 16'h200;
			16'h4ca4: y = 16'h200;
			16'h4ca5: y = 16'h200;
			16'h4ca6: y = 16'h200;
			16'h4ca7: y = 16'h200;
			16'h4ca8: y = 16'h200;
			16'h4ca9: y = 16'h200;
			16'h4caa: y = 16'h200;
			16'h4cab: y = 16'h200;
			16'h4cac: y = 16'h200;
			16'h4cad: y = 16'h200;
			16'h4cae: y = 16'h200;
			16'h4caf: y = 16'h200;
			16'h4cb0: y = 16'h200;
			16'h4cb1: y = 16'h200;
			16'h4cb2: y = 16'h200;
			16'h4cb3: y = 16'h200;
			16'h4cb4: y = 16'h200;
			16'h4cb5: y = 16'h200;
			16'h4cb6: y = 16'h200;
			16'h4cb7: y = 16'h200;
			16'h4cb8: y = 16'h200;
			16'h4cb9: y = 16'h200;
			16'h4cba: y = 16'h200;
			16'h4cbb: y = 16'h200;
			16'h4cbc: y = 16'h200;
			16'h4cbd: y = 16'h200;
			16'h4cbe: y = 16'h200;
			16'h4cbf: y = 16'h200;
			16'h4cc0: y = 16'h200;
			16'h4cc1: y = 16'h200;
			16'h4cc2: y = 16'h200;
			16'h4cc3: y = 16'h200;
			16'h4cc4: y = 16'h200;
			16'h4cc5: y = 16'h200;
			16'h4cc6: y = 16'h200;
			16'h4cc7: y = 16'h200;
			16'h4cc8: y = 16'h200;
			16'h4cc9: y = 16'h200;
			16'h4cca: y = 16'h200;
			16'h4ccb: y = 16'h200;
			16'h4ccc: y = 16'h200;
			16'h4ccd: y = 16'h200;
			16'h4cce: y = 16'h200;
			16'h4ccf: y = 16'h200;
			16'h4cd0: y = 16'h200;
			16'h4cd1: y = 16'h200;
			16'h4cd2: y = 16'h200;
			16'h4cd3: y = 16'h200;
			16'h4cd4: y = 16'h200;
			16'h4cd5: y = 16'h200;
			16'h4cd6: y = 16'h200;
			16'h4cd7: y = 16'h200;
			16'h4cd8: y = 16'h200;
			16'h4cd9: y = 16'h200;
			16'h4cda: y = 16'h200;
			16'h4cdb: y = 16'h200;
			16'h4cdc: y = 16'h200;
			16'h4cdd: y = 16'h200;
			16'h4cde: y = 16'h200;
			16'h4cdf: y = 16'h200;
			16'h4ce0: y = 16'h200;
			16'h4ce1: y = 16'h200;
			16'h4ce2: y = 16'h200;
			16'h4ce3: y = 16'h200;
			16'h4ce4: y = 16'h200;
			16'h4ce5: y = 16'h200;
			16'h4ce6: y = 16'h200;
			16'h4ce7: y = 16'h200;
			16'h4ce8: y = 16'h200;
			16'h4ce9: y = 16'h200;
			16'h4cea: y = 16'h200;
			16'h4ceb: y = 16'h200;
			16'h4cec: y = 16'h200;
			16'h4ced: y = 16'h200;
			16'h4cee: y = 16'h200;
			16'h4cef: y = 16'h200;
			16'h4cf0: y = 16'h200;
			16'h4cf1: y = 16'h200;
			16'h4cf2: y = 16'h200;
			16'h4cf3: y = 16'h200;
			16'h4cf4: y = 16'h200;
			16'h4cf5: y = 16'h200;
			16'h4cf6: y = 16'h200;
			16'h4cf7: y = 16'h200;
			16'h4cf8: y = 16'h200;
			16'h4cf9: y = 16'h200;
			16'h4cfa: y = 16'h200;
			16'h4cfb: y = 16'h200;
			16'h4cfc: y = 16'h200;
			16'h4cfd: y = 16'h200;
			16'h4cfe: y = 16'h200;
			16'h4cff: y = 16'h200;
			16'h4d00: y = 16'h200;
			16'h4d01: y = 16'h200;
			16'h4d02: y = 16'h200;
			16'h4d03: y = 16'h200;
			16'h4d04: y = 16'h200;
			16'h4d05: y = 16'h200;
			16'h4d06: y = 16'h200;
			16'h4d07: y = 16'h200;
			16'h4d08: y = 16'h200;
			16'h4d09: y = 16'h200;
			16'h4d0a: y = 16'h200;
			16'h4d0b: y = 16'h200;
			16'h4d0c: y = 16'h200;
			16'h4d0d: y = 16'h200;
			16'h4d0e: y = 16'h200;
			16'h4d0f: y = 16'h200;
			16'h4d10: y = 16'h200;
			16'h4d11: y = 16'h200;
			16'h4d12: y = 16'h200;
			16'h4d13: y = 16'h200;
			16'h4d14: y = 16'h200;
			16'h4d15: y = 16'h200;
			16'h4d16: y = 16'h200;
			16'h4d17: y = 16'h200;
			16'h4d18: y = 16'h200;
			16'h4d19: y = 16'h200;
			16'h4d1a: y = 16'h200;
			16'h4d1b: y = 16'h200;
			16'h4d1c: y = 16'h200;
			16'h4d1d: y = 16'h200;
			16'h4d1e: y = 16'h200;
			16'h4d1f: y = 16'h200;
			16'h4d20: y = 16'h200;
			16'h4d21: y = 16'h200;
			16'h4d22: y = 16'h200;
			16'h4d23: y = 16'h200;
			16'h4d24: y = 16'h200;
			16'h4d25: y = 16'h200;
			16'h4d26: y = 16'h200;
			16'h4d27: y = 16'h200;
			16'h4d28: y = 16'h200;
			16'h4d29: y = 16'h200;
			16'h4d2a: y = 16'h200;
			16'h4d2b: y = 16'h200;
			16'h4d2c: y = 16'h200;
			16'h4d2d: y = 16'h200;
			16'h4d2e: y = 16'h200;
			16'h4d2f: y = 16'h200;
			16'h4d30: y = 16'h200;
			16'h4d31: y = 16'h200;
			16'h4d32: y = 16'h200;
			16'h4d33: y = 16'h200;
			16'h4d34: y = 16'h200;
			16'h4d35: y = 16'h200;
			16'h4d36: y = 16'h200;
			16'h4d37: y = 16'h200;
			16'h4d38: y = 16'h200;
			16'h4d39: y = 16'h200;
			16'h4d3a: y = 16'h200;
			16'h4d3b: y = 16'h200;
			16'h4d3c: y = 16'h200;
			16'h4d3d: y = 16'h200;
			16'h4d3e: y = 16'h200;
			16'h4d3f: y = 16'h200;
			16'h4d40: y = 16'h200;
			16'h4d41: y = 16'h200;
			16'h4d42: y = 16'h200;
			16'h4d43: y = 16'h200;
			16'h4d44: y = 16'h200;
			16'h4d45: y = 16'h200;
			16'h4d46: y = 16'h200;
			16'h4d47: y = 16'h200;
			16'h4d48: y = 16'h200;
			16'h4d49: y = 16'h200;
			16'h4d4a: y = 16'h200;
			16'h4d4b: y = 16'h200;
			16'h4d4c: y = 16'h200;
			16'h4d4d: y = 16'h200;
			16'h4d4e: y = 16'h200;
			16'h4d4f: y = 16'h200;
			16'h4d50: y = 16'h200;
			16'h4d51: y = 16'h200;
			16'h4d52: y = 16'h200;
			16'h4d53: y = 16'h200;
			16'h4d54: y = 16'h200;
			16'h4d55: y = 16'h200;
			16'h4d56: y = 16'h200;
			16'h4d57: y = 16'h200;
			16'h4d58: y = 16'h200;
			16'h4d59: y = 16'h200;
			16'h4d5a: y = 16'h200;
			16'h4d5b: y = 16'h200;
			16'h4d5c: y = 16'h200;
			16'h4d5d: y = 16'h200;
			16'h4d5e: y = 16'h200;
			16'h4d5f: y = 16'h200;
			16'h4d60: y = 16'h200;
			16'h4d61: y = 16'h200;
			16'h4d62: y = 16'h200;
			16'h4d63: y = 16'h200;
			16'h4d64: y = 16'h200;
			16'h4d65: y = 16'h200;
			16'h4d66: y = 16'h200;
			16'h4d67: y = 16'h200;
			16'h4d68: y = 16'h200;
			16'h4d69: y = 16'h200;
			16'h4d6a: y = 16'h200;
			16'h4d6b: y = 16'h200;
			16'h4d6c: y = 16'h200;
			16'h4d6d: y = 16'h200;
			16'h4d6e: y = 16'h200;
			16'h4d6f: y = 16'h200;
			16'h4d70: y = 16'h200;
			16'h4d71: y = 16'h200;
			16'h4d72: y = 16'h200;
			16'h4d73: y = 16'h200;
			16'h4d74: y = 16'h200;
			16'h4d75: y = 16'h200;
			16'h4d76: y = 16'h200;
			16'h4d77: y = 16'h200;
			16'h4d78: y = 16'h200;
			16'h4d79: y = 16'h200;
			16'h4d7a: y = 16'h200;
			16'h4d7b: y = 16'h200;
			16'h4d7c: y = 16'h200;
			16'h4d7d: y = 16'h200;
			16'h4d7e: y = 16'h200;
			16'h4d7f: y = 16'h200;
			16'h4d80: y = 16'h200;
			16'h4d81: y = 16'h200;
			16'h4d82: y = 16'h200;
			16'h4d83: y = 16'h200;
			16'h4d84: y = 16'h200;
			16'h4d85: y = 16'h200;
			16'h4d86: y = 16'h200;
			16'h4d87: y = 16'h200;
			16'h4d88: y = 16'h200;
			16'h4d89: y = 16'h200;
			16'h4d8a: y = 16'h200;
			16'h4d8b: y = 16'h200;
			16'h4d8c: y = 16'h200;
			16'h4d8d: y = 16'h200;
			16'h4d8e: y = 16'h200;
			16'h4d8f: y = 16'h200;
			16'h4d90: y = 16'h200;
			16'h4d91: y = 16'h200;
			16'h4d92: y = 16'h200;
			16'h4d93: y = 16'h200;
			16'h4d94: y = 16'h200;
			16'h4d95: y = 16'h200;
			16'h4d96: y = 16'h200;
			16'h4d97: y = 16'h200;
			16'h4d98: y = 16'h200;
			16'h4d99: y = 16'h200;
			16'h4d9a: y = 16'h200;
			16'h4d9b: y = 16'h200;
			16'h4d9c: y = 16'h200;
			16'h4d9d: y = 16'h200;
			16'h4d9e: y = 16'h200;
			16'h4d9f: y = 16'h200;
			16'h4da0: y = 16'h200;
			16'h4da1: y = 16'h200;
			16'h4da2: y = 16'h200;
			16'h4da3: y = 16'h200;
			16'h4da4: y = 16'h200;
			16'h4da5: y = 16'h200;
			16'h4da6: y = 16'h200;
			16'h4da7: y = 16'h200;
			16'h4da8: y = 16'h200;
			16'h4da9: y = 16'h200;
			16'h4daa: y = 16'h200;
			16'h4dab: y = 16'h200;
			16'h4dac: y = 16'h200;
			16'h4dad: y = 16'h200;
			16'h4dae: y = 16'h200;
			16'h4daf: y = 16'h200;
			16'h4db0: y = 16'h200;
			16'h4db1: y = 16'h200;
			16'h4db2: y = 16'h200;
			16'h4db3: y = 16'h200;
			16'h4db4: y = 16'h200;
			16'h4db5: y = 16'h200;
			16'h4db6: y = 16'h200;
			16'h4db7: y = 16'h200;
			16'h4db8: y = 16'h200;
			16'h4db9: y = 16'h200;
			16'h4dba: y = 16'h200;
			16'h4dbb: y = 16'h200;
			16'h4dbc: y = 16'h200;
			16'h4dbd: y = 16'h200;
			16'h4dbe: y = 16'h200;
			16'h4dbf: y = 16'h200;
			16'h4dc0: y = 16'h200;
			16'h4dc1: y = 16'h200;
			16'h4dc2: y = 16'h200;
			16'h4dc3: y = 16'h200;
			16'h4dc4: y = 16'h200;
			16'h4dc5: y = 16'h200;
			16'h4dc6: y = 16'h200;
			16'h4dc7: y = 16'h200;
			16'h4dc8: y = 16'h200;
			16'h4dc9: y = 16'h200;
			16'h4dca: y = 16'h200;
			16'h4dcb: y = 16'h200;
			16'h4dcc: y = 16'h200;
			16'h4dcd: y = 16'h200;
			16'h4dce: y = 16'h200;
			16'h4dcf: y = 16'h200;
			16'h4dd0: y = 16'h200;
			16'h4dd1: y = 16'h200;
			16'h4dd2: y = 16'h200;
			16'h4dd3: y = 16'h200;
			16'h4dd4: y = 16'h200;
			16'h4dd5: y = 16'h200;
			16'h4dd6: y = 16'h200;
			16'h4dd7: y = 16'h200;
			16'h4dd8: y = 16'h200;
			16'h4dd9: y = 16'h200;
			16'h4dda: y = 16'h200;
			16'h4ddb: y = 16'h200;
			16'h4ddc: y = 16'h200;
			16'h4ddd: y = 16'h200;
			16'h4dde: y = 16'h200;
			16'h4ddf: y = 16'h200;
			16'h4de0: y = 16'h200;
			16'h4de1: y = 16'h200;
			16'h4de2: y = 16'h200;
			16'h4de3: y = 16'h200;
			16'h4de4: y = 16'h200;
			16'h4de5: y = 16'h200;
			16'h4de6: y = 16'h200;
			16'h4de7: y = 16'h200;
			16'h4de8: y = 16'h200;
			16'h4de9: y = 16'h200;
			16'h4dea: y = 16'h200;
			16'h4deb: y = 16'h200;
			16'h4dec: y = 16'h200;
			16'h4ded: y = 16'h200;
			16'h4dee: y = 16'h200;
			16'h4def: y = 16'h200;
			16'h4df0: y = 16'h200;
			16'h4df1: y = 16'h200;
			16'h4df2: y = 16'h200;
			16'h4df3: y = 16'h200;
			16'h4df4: y = 16'h200;
			16'h4df5: y = 16'h200;
			16'h4df6: y = 16'h200;
			16'h4df7: y = 16'h200;
			16'h4df8: y = 16'h200;
			16'h4df9: y = 16'h200;
			16'h4dfa: y = 16'h200;
			16'h4dfb: y = 16'h200;
			16'h4dfc: y = 16'h200;
			16'h4dfd: y = 16'h200;
			16'h4dfe: y = 16'h200;
			16'h4dff: y = 16'h200;
			16'h4e00: y = 16'h200;
			16'h4e01: y = 16'h200;
			16'h4e02: y = 16'h200;
			16'h4e03: y = 16'h200;
			16'h4e04: y = 16'h200;
			16'h4e05: y = 16'h200;
			16'h4e06: y = 16'h200;
			16'h4e07: y = 16'h200;
			16'h4e08: y = 16'h200;
			16'h4e09: y = 16'h200;
			16'h4e0a: y = 16'h200;
			16'h4e0b: y = 16'h200;
			16'h4e0c: y = 16'h200;
			16'h4e0d: y = 16'h200;
			16'h4e0e: y = 16'h200;
			16'h4e0f: y = 16'h200;
			16'h4e10: y = 16'h200;
			16'h4e11: y = 16'h200;
			16'h4e12: y = 16'h200;
			16'h4e13: y = 16'h200;
			16'h4e14: y = 16'h200;
			16'h4e15: y = 16'h200;
			16'h4e16: y = 16'h200;
			16'h4e17: y = 16'h200;
			16'h4e18: y = 16'h200;
			16'h4e19: y = 16'h200;
			16'h4e1a: y = 16'h200;
			16'h4e1b: y = 16'h200;
			16'h4e1c: y = 16'h200;
			16'h4e1d: y = 16'h200;
			16'h4e1e: y = 16'h200;
			16'h4e1f: y = 16'h200;
			16'h4e20: y = 16'h200;
			16'h4e21: y = 16'h200;
			16'h4e22: y = 16'h200;
			16'h4e23: y = 16'h200;
			16'h4e24: y = 16'h200;
			16'h4e25: y = 16'h200;
			16'h4e26: y = 16'h200;
			16'h4e27: y = 16'h200;
			16'h4e28: y = 16'h200;
			16'h4e29: y = 16'h200;
			16'h4e2a: y = 16'h200;
			16'h4e2b: y = 16'h200;
			16'h4e2c: y = 16'h200;
			16'h4e2d: y = 16'h200;
			16'h4e2e: y = 16'h200;
			16'h4e2f: y = 16'h200;
			16'h4e30: y = 16'h200;
			16'h4e31: y = 16'h200;
			16'h4e32: y = 16'h200;
			16'h4e33: y = 16'h200;
			16'h4e34: y = 16'h200;
			16'h4e35: y = 16'h200;
			16'h4e36: y = 16'h200;
			16'h4e37: y = 16'h200;
			16'h4e38: y = 16'h200;
			16'h4e39: y = 16'h200;
			16'h4e3a: y = 16'h200;
			16'h4e3b: y = 16'h200;
			16'h4e3c: y = 16'h200;
			16'h4e3d: y = 16'h200;
			16'h4e3e: y = 16'h200;
			16'h4e3f: y = 16'h200;
			16'h4e40: y = 16'h200;
			16'h4e41: y = 16'h200;
			16'h4e42: y = 16'h200;
			16'h4e43: y = 16'h200;
			16'h4e44: y = 16'h200;
			16'h4e45: y = 16'h200;
			16'h4e46: y = 16'h200;
			16'h4e47: y = 16'h200;
			16'h4e48: y = 16'h200;
			16'h4e49: y = 16'h200;
			16'h4e4a: y = 16'h200;
			16'h4e4b: y = 16'h200;
			16'h4e4c: y = 16'h200;
			16'h4e4d: y = 16'h200;
			16'h4e4e: y = 16'h200;
			16'h4e4f: y = 16'h200;
			16'h4e50: y = 16'h200;
			16'h4e51: y = 16'h200;
			16'h4e52: y = 16'h200;
			16'h4e53: y = 16'h200;
			16'h4e54: y = 16'h200;
			16'h4e55: y = 16'h200;
			16'h4e56: y = 16'h200;
			16'h4e57: y = 16'h200;
			16'h4e58: y = 16'h200;
			16'h4e59: y = 16'h200;
			16'h4e5a: y = 16'h200;
			16'h4e5b: y = 16'h200;
			16'h4e5c: y = 16'h200;
			16'h4e5d: y = 16'h200;
			16'h4e5e: y = 16'h200;
			16'h4e5f: y = 16'h200;
			16'h4e60: y = 16'h200;
			16'h4e61: y = 16'h200;
			16'h4e62: y = 16'h200;
			16'h4e63: y = 16'h200;
			16'h4e64: y = 16'h200;
			16'h4e65: y = 16'h200;
			16'h4e66: y = 16'h200;
			16'h4e67: y = 16'h200;
			16'h4e68: y = 16'h200;
			16'h4e69: y = 16'h200;
			16'h4e6a: y = 16'h200;
			16'h4e6b: y = 16'h200;
			16'h4e6c: y = 16'h200;
			16'h4e6d: y = 16'h200;
			16'h4e6e: y = 16'h200;
			16'h4e6f: y = 16'h200;
			16'h4e70: y = 16'h200;
			16'h4e71: y = 16'h200;
			16'h4e72: y = 16'h200;
			16'h4e73: y = 16'h200;
			16'h4e74: y = 16'h200;
			16'h4e75: y = 16'h200;
			16'h4e76: y = 16'h200;
			16'h4e77: y = 16'h200;
			16'h4e78: y = 16'h200;
			16'h4e79: y = 16'h200;
			16'h4e7a: y = 16'h200;
			16'h4e7b: y = 16'h200;
			16'h4e7c: y = 16'h200;
			16'h4e7d: y = 16'h200;
			16'h4e7e: y = 16'h200;
			16'h4e7f: y = 16'h200;
			16'h4e80: y = 16'h200;
			16'h4e81: y = 16'h200;
			16'h4e82: y = 16'h200;
			16'h4e83: y = 16'h200;
			16'h4e84: y = 16'h200;
			16'h4e85: y = 16'h200;
			16'h4e86: y = 16'h200;
			16'h4e87: y = 16'h200;
			16'h4e88: y = 16'h200;
			16'h4e89: y = 16'h200;
			16'h4e8a: y = 16'h200;
			16'h4e8b: y = 16'h200;
			16'h4e8c: y = 16'h200;
			16'h4e8d: y = 16'h200;
			16'h4e8e: y = 16'h200;
			16'h4e8f: y = 16'h200;
			16'h4e90: y = 16'h200;
			16'h4e91: y = 16'h200;
			16'h4e92: y = 16'h200;
			16'h4e93: y = 16'h200;
			16'h4e94: y = 16'h200;
			16'h4e95: y = 16'h200;
			16'h4e96: y = 16'h200;
			16'h4e97: y = 16'h200;
			16'h4e98: y = 16'h200;
			16'h4e99: y = 16'h200;
			16'h4e9a: y = 16'h200;
			16'h4e9b: y = 16'h200;
			16'h4e9c: y = 16'h200;
			16'h4e9d: y = 16'h200;
			16'h4e9e: y = 16'h200;
			16'h4e9f: y = 16'h200;
			16'h4ea0: y = 16'h200;
			16'h4ea1: y = 16'h200;
			16'h4ea2: y = 16'h200;
			16'h4ea3: y = 16'h200;
			16'h4ea4: y = 16'h200;
			16'h4ea5: y = 16'h200;
			16'h4ea6: y = 16'h200;
			16'h4ea7: y = 16'h200;
			16'h4ea8: y = 16'h200;
			16'h4ea9: y = 16'h200;
			16'h4eaa: y = 16'h200;
			16'h4eab: y = 16'h200;
			16'h4eac: y = 16'h200;
			16'h4ead: y = 16'h200;
			16'h4eae: y = 16'h200;
			16'h4eaf: y = 16'h200;
			16'h4eb0: y = 16'h200;
			16'h4eb1: y = 16'h200;
			16'h4eb2: y = 16'h200;
			16'h4eb3: y = 16'h200;
			16'h4eb4: y = 16'h200;
			16'h4eb5: y = 16'h200;
			16'h4eb6: y = 16'h200;
			16'h4eb7: y = 16'h200;
			16'h4eb8: y = 16'h200;
			16'h4eb9: y = 16'h200;
			16'h4eba: y = 16'h200;
			16'h4ebb: y = 16'h200;
			16'h4ebc: y = 16'h200;
			16'h4ebd: y = 16'h200;
			16'h4ebe: y = 16'h200;
			16'h4ebf: y = 16'h200;
			16'h4ec0: y = 16'h200;
			16'h4ec1: y = 16'h200;
			16'h4ec2: y = 16'h200;
			16'h4ec3: y = 16'h200;
			16'h4ec4: y = 16'h200;
			16'h4ec5: y = 16'h200;
			16'h4ec6: y = 16'h200;
			16'h4ec7: y = 16'h200;
			16'h4ec8: y = 16'h200;
			16'h4ec9: y = 16'h200;
			16'h4eca: y = 16'h200;
			16'h4ecb: y = 16'h200;
			16'h4ecc: y = 16'h200;
			16'h4ecd: y = 16'h200;
			16'h4ece: y = 16'h200;
			16'h4ecf: y = 16'h200;
			16'h4ed0: y = 16'h200;
			16'h4ed1: y = 16'h200;
			16'h4ed2: y = 16'h200;
			16'h4ed3: y = 16'h200;
			16'h4ed4: y = 16'h200;
			16'h4ed5: y = 16'h200;
			16'h4ed6: y = 16'h200;
			16'h4ed7: y = 16'h200;
			16'h4ed8: y = 16'h200;
			16'h4ed9: y = 16'h200;
			16'h4eda: y = 16'h200;
			16'h4edb: y = 16'h200;
			16'h4edc: y = 16'h200;
			16'h4edd: y = 16'h200;
			16'h4ede: y = 16'h200;
			16'h4edf: y = 16'h200;
			16'h4ee0: y = 16'h200;
			16'h4ee1: y = 16'h200;
			16'h4ee2: y = 16'h200;
			16'h4ee3: y = 16'h200;
			16'h4ee4: y = 16'h200;
			16'h4ee5: y = 16'h200;
			16'h4ee6: y = 16'h200;
			16'h4ee7: y = 16'h200;
			16'h4ee8: y = 16'h200;
			16'h4ee9: y = 16'h200;
			16'h4eea: y = 16'h200;
			16'h4eeb: y = 16'h200;
			16'h4eec: y = 16'h200;
			16'h4eed: y = 16'h200;
			16'h4eee: y = 16'h200;
			16'h4eef: y = 16'h200;
			16'h4ef0: y = 16'h200;
			16'h4ef1: y = 16'h200;
			16'h4ef2: y = 16'h200;
			16'h4ef3: y = 16'h200;
			16'h4ef4: y = 16'h200;
			16'h4ef5: y = 16'h200;
			16'h4ef6: y = 16'h200;
			16'h4ef7: y = 16'h200;
			16'h4ef8: y = 16'h200;
			16'h4ef9: y = 16'h200;
			16'h4efa: y = 16'h200;
			16'h4efb: y = 16'h200;
			16'h4efc: y = 16'h200;
			16'h4efd: y = 16'h200;
			16'h4efe: y = 16'h200;
			16'h4eff: y = 16'h200;
			16'h4f00: y = 16'h200;
			16'h4f01: y = 16'h200;
			16'h4f02: y = 16'h200;
			16'h4f03: y = 16'h200;
			16'h4f04: y = 16'h200;
			16'h4f05: y = 16'h200;
			16'h4f06: y = 16'h200;
			16'h4f07: y = 16'h200;
			16'h4f08: y = 16'h200;
			16'h4f09: y = 16'h200;
			16'h4f0a: y = 16'h200;
			16'h4f0b: y = 16'h200;
			16'h4f0c: y = 16'h200;
			16'h4f0d: y = 16'h200;
			16'h4f0e: y = 16'h200;
			16'h4f0f: y = 16'h200;
			16'h4f10: y = 16'h200;
			16'h4f11: y = 16'h200;
			16'h4f12: y = 16'h200;
			16'h4f13: y = 16'h200;
			16'h4f14: y = 16'h200;
			16'h4f15: y = 16'h200;
			16'h4f16: y = 16'h200;
			16'h4f17: y = 16'h200;
			16'h4f18: y = 16'h200;
			16'h4f19: y = 16'h200;
			16'h4f1a: y = 16'h200;
			16'h4f1b: y = 16'h200;
			16'h4f1c: y = 16'h200;
			16'h4f1d: y = 16'h200;
			16'h4f1e: y = 16'h200;
			16'h4f1f: y = 16'h200;
			16'h4f20: y = 16'h200;
			16'h4f21: y = 16'h200;
			16'h4f22: y = 16'h200;
			16'h4f23: y = 16'h200;
			16'h4f24: y = 16'h200;
			16'h4f25: y = 16'h200;
			16'h4f26: y = 16'h200;
			16'h4f27: y = 16'h200;
			16'h4f28: y = 16'h200;
			16'h4f29: y = 16'h200;
			16'h4f2a: y = 16'h200;
			16'h4f2b: y = 16'h200;
			16'h4f2c: y = 16'h200;
			16'h4f2d: y = 16'h200;
			16'h4f2e: y = 16'h200;
			16'h4f2f: y = 16'h200;
			16'h4f30: y = 16'h200;
			16'h4f31: y = 16'h200;
			16'h4f32: y = 16'h200;
			16'h4f33: y = 16'h200;
			16'h4f34: y = 16'h200;
			16'h4f35: y = 16'h200;
			16'h4f36: y = 16'h200;
			16'h4f37: y = 16'h200;
			16'h4f38: y = 16'h200;
			16'h4f39: y = 16'h200;
			16'h4f3a: y = 16'h200;
			16'h4f3b: y = 16'h200;
			16'h4f3c: y = 16'h200;
			16'h4f3d: y = 16'h200;
			16'h4f3e: y = 16'h200;
			16'h4f3f: y = 16'h200;
			16'h4f40: y = 16'h200;
			16'h4f41: y = 16'h200;
			16'h4f42: y = 16'h200;
			16'h4f43: y = 16'h200;
			16'h4f44: y = 16'h200;
			16'h4f45: y = 16'h200;
			16'h4f46: y = 16'h200;
			16'h4f47: y = 16'h200;
			16'h4f48: y = 16'h200;
			16'h4f49: y = 16'h200;
			16'h4f4a: y = 16'h200;
			16'h4f4b: y = 16'h200;
			16'h4f4c: y = 16'h200;
			16'h4f4d: y = 16'h200;
			16'h4f4e: y = 16'h200;
			16'h4f4f: y = 16'h200;
			16'h4f50: y = 16'h200;
			16'h4f51: y = 16'h200;
			16'h4f52: y = 16'h200;
			16'h4f53: y = 16'h200;
			16'h4f54: y = 16'h200;
			16'h4f55: y = 16'h200;
			16'h4f56: y = 16'h200;
			16'h4f57: y = 16'h200;
			16'h4f58: y = 16'h200;
			16'h4f59: y = 16'h200;
			16'h4f5a: y = 16'h200;
			16'h4f5b: y = 16'h200;
			16'h4f5c: y = 16'h200;
			16'h4f5d: y = 16'h200;
			16'h4f5e: y = 16'h200;
			16'h4f5f: y = 16'h200;
			16'h4f60: y = 16'h200;
			16'h4f61: y = 16'h200;
			16'h4f62: y = 16'h200;
			16'h4f63: y = 16'h200;
			16'h4f64: y = 16'h200;
			16'h4f65: y = 16'h200;
			16'h4f66: y = 16'h200;
			16'h4f67: y = 16'h200;
			16'h4f68: y = 16'h200;
			16'h4f69: y = 16'h200;
			16'h4f6a: y = 16'h200;
			16'h4f6b: y = 16'h200;
			16'h4f6c: y = 16'h200;
			16'h4f6d: y = 16'h200;
			16'h4f6e: y = 16'h200;
			16'h4f6f: y = 16'h200;
			16'h4f70: y = 16'h200;
			16'h4f71: y = 16'h200;
			16'h4f72: y = 16'h200;
			16'h4f73: y = 16'h200;
			16'h4f74: y = 16'h200;
			16'h4f75: y = 16'h200;
			16'h4f76: y = 16'h200;
			16'h4f77: y = 16'h200;
			16'h4f78: y = 16'h200;
			16'h4f79: y = 16'h200;
			16'h4f7a: y = 16'h200;
			16'h4f7b: y = 16'h200;
			16'h4f7c: y = 16'h200;
			16'h4f7d: y = 16'h200;
			16'h4f7e: y = 16'h200;
			16'h4f7f: y = 16'h200;
			16'h4f80: y = 16'h200;
			16'h4f81: y = 16'h200;
			16'h4f82: y = 16'h200;
			16'h4f83: y = 16'h200;
			16'h4f84: y = 16'h200;
			16'h4f85: y = 16'h200;
			16'h4f86: y = 16'h200;
			16'h4f87: y = 16'h200;
			16'h4f88: y = 16'h200;
			16'h4f89: y = 16'h200;
			16'h4f8a: y = 16'h200;
			16'h4f8b: y = 16'h200;
			16'h4f8c: y = 16'h200;
			16'h4f8d: y = 16'h200;
			16'h4f8e: y = 16'h200;
			16'h4f8f: y = 16'h200;
			16'h4f90: y = 16'h200;
			16'h4f91: y = 16'h200;
			16'h4f92: y = 16'h200;
			16'h4f93: y = 16'h200;
			16'h4f94: y = 16'h200;
			16'h4f95: y = 16'h200;
			16'h4f96: y = 16'h200;
			16'h4f97: y = 16'h200;
			16'h4f98: y = 16'h200;
			16'h4f99: y = 16'h200;
			16'h4f9a: y = 16'h200;
			16'h4f9b: y = 16'h200;
			16'h4f9c: y = 16'h200;
			16'h4f9d: y = 16'h200;
			16'h4f9e: y = 16'h200;
			16'h4f9f: y = 16'h200;
			16'h4fa0: y = 16'h200;
			16'h4fa1: y = 16'h200;
			16'h4fa2: y = 16'h200;
			16'h4fa3: y = 16'h200;
			16'h4fa4: y = 16'h200;
			16'h4fa5: y = 16'h200;
			16'h4fa6: y = 16'h200;
			16'h4fa7: y = 16'h200;
			16'h4fa8: y = 16'h200;
			16'h4fa9: y = 16'h200;
			16'h4faa: y = 16'h200;
			16'h4fab: y = 16'h200;
			16'h4fac: y = 16'h200;
			16'h4fad: y = 16'h200;
			16'h4fae: y = 16'h200;
			16'h4faf: y = 16'h200;
			16'h4fb0: y = 16'h200;
			16'h4fb1: y = 16'h200;
			16'h4fb2: y = 16'h200;
			16'h4fb3: y = 16'h200;
			16'h4fb4: y = 16'h200;
			16'h4fb5: y = 16'h200;
			16'h4fb6: y = 16'h200;
			16'h4fb7: y = 16'h200;
			16'h4fb8: y = 16'h200;
			16'h4fb9: y = 16'h200;
			16'h4fba: y = 16'h200;
			16'h4fbb: y = 16'h200;
			16'h4fbc: y = 16'h200;
			16'h4fbd: y = 16'h200;
			16'h4fbe: y = 16'h200;
			16'h4fbf: y = 16'h200;
			16'h4fc0: y = 16'h200;
			16'h4fc1: y = 16'h200;
			16'h4fc2: y = 16'h200;
			16'h4fc3: y = 16'h200;
			16'h4fc4: y = 16'h200;
			16'h4fc5: y = 16'h200;
			16'h4fc6: y = 16'h200;
			16'h4fc7: y = 16'h200;
			16'h4fc8: y = 16'h200;
			16'h4fc9: y = 16'h200;
			16'h4fca: y = 16'h200;
			16'h4fcb: y = 16'h200;
			16'h4fcc: y = 16'h200;
			16'h4fcd: y = 16'h200;
			16'h4fce: y = 16'h200;
			16'h4fcf: y = 16'h200;
			16'h4fd0: y = 16'h200;
			16'h4fd1: y = 16'h200;
			16'h4fd2: y = 16'h200;
			16'h4fd3: y = 16'h200;
			16'h4fd4: y = 16'h200;
			16'h4fd5: y = 16'h200;
			16'h4fd6: y = 16'h200;
			16'h4fd7: y = 16'h200;
			16'h4fd8: y = 16'h200;
			16'h4fd9: y = 16'h200;
			16'h4fda: y = 16'h200;
			16'h4fdb: y = 16'h200;
			16'h4fdc: y = 16'h200;
			16'h4fdd: y = 16'h200;
			16'h4fde: y = 16'h200;
			16'h4fdf: y = 16'h200;
			16'h4fe0: y = 16'h200;
			16'h4fe1: y = 16'h200;
			16'h4fe2: y = 16'h200;
			16'h4fe3: y = 16'h200;
			16'h4fe4: y = 16'h200;
			16'h4fe5: y = 16'h200;
			16'h4fe6: y = 16'h200;
			16'h4fe7: y = 16'h200;
			16'h4fe8: y = 16'h200;
			16'h4fe9: y = 16'h200;
			16'h4fea: y = 16'h200;
			16'h4feb: y = 16'h200;
			16'h4fec: y = 16'h200;
			16'h4fed: y = 16'h200;
			16'h4fee: y = 16'h200;
			16'h4fef: y = 16'h200;
			16'h4ff0: y = 16'h200;
			16'h4ff1: y = 16'h200;
			16'h4ff2: y = 16'h200;
			16'h4ff3: y = 16'h200;
			16'h4ff4: y = 16'h200;
			16'h4ff5: y = 16'h200;
			16'h4ff6: y = 16'h200;
			16'h4ff7: y = 16'h200;
			16'h4ff8: y = 16'h200;
			16'h4ff9: y = 16'h200;
			16'h4ffa: y = 16'h200;
			16'h4ffb: y = 16'h200;
			16'h4ffc: y = 16'h200;
			16'h4ffd: y = 16'h200;
			16'h4ffe: y = 16'h200;
			16'h4fff: y = 16'h200;
			16'h5000: y = 16'h200;
			16'h5001: y = 16'h200;
			16'h5002: y = 16'h200;
			16'h5003: y = 16'h200;
			16'h5004: y = 16'h200;
			16'h5005: y = 16'h200;
			16'h5006: y = 16'h200;
			16'h5007: y = 16'h200;
			16'h5008: y = 16'h200;
			16'h5009: y = 16'h200;
			16'h500a: y = 16'h200;
			16'h500b: y = 16'h200;
			16'h500c: y = 16'h200;
			16'h500d: y = 16'h200;
			16'h500e: y = 16'h200;
			16'h500f: y = 16'h200;
			16'h5010: y = 16'h200;
			16'h5011: y = 16'h200;
			16'h5012: y = 16'h200;
			16'h5013: y = 16'h200;
			16'h5014: y = 16'h200;
			16'h5015: y = 16'h200;
			16'h5016: y = 16'h200;
			16'h5017: y = 16'h200;
			16'h5018: y = 16'h200;
			16'h5019: y = 16'h200;
			16'h501a: y = 16'h200;
			16'h501b: y = 16'h200;
			16'h501c: y = 16'h200;
			16'h501d: y = 16'h200;
			16'h501e: y = 16'h200;
			16'h501f: y = 16'h200;
			16'h5020: y = 16'h200;
			16'h5021: y = 16'h200;
			16'h5022: y = 16'h200;
			16'h5023: y = 16'h200;
			16'h5024: y = 16'h200;
			16'h5025: y = 16'h200;
			16'h5026: y = 16'h200;
			16'h5027: y = 16'h200;
			16'h5028: y = 16'h200;
			16'h5029: y = 16'h200;
			16'h502a: y = 16'h200;
			16'h502b: y = 16'h200;
			16'h502c: y = 16'h200;
			16'h502d: y = 16'h200;
			16'h502e: y = 16'h200;
			16'h502f: y = 16'h200;
			16'h5030: y = 16'h200;
			16'h5031: y = 16'h200;
			16'h5032: y = 16'h200;
			16'h5033: y = 16'h200;
			16'h5034: y = 16'h200;
			16'h5035: y = 16'h200;
			16'h5036: y = 16'h200;
			16'h5037: y = 16'h200;
			16'h5038: y = 16'h200;
			16'h5039: y = 16'h200;
			16'h503a: y = 16'h200;
			16'h503b: y = 16'h200;
			16'h503c: y = 16'h200;
			16'h503d: y = 16'h200;
			16'h503e: y = 16'h200;
			16'h503f: y = 16'h200;
			16'h5040: y = 16'h200;
			16'h5041: y = 16'h200;
			16'h5042: y = 16'h200;
			16'h5043: y = 16'h200;
			16'h5044: y = 16'h200;
			16'h5045: y = 16'h200;
			16'h5046: y = 16'h200;
			16'h5047: y = 16'h200;
			16'h5048: y = 16'h200;
			16'h5049: y = 16'h200;
			16'h504a: y = 16'h200;
			16'h504b: y = 16'h200;
			16'h504c: y = 16'h200;
			16'h504d: y = 16'h200;
			16'h504e: y = 16'h200;
			16'h504f: y = 16'h200;
			16'h5050: y = 16'h200;
			16'h5051: y = 16'h200;
			16'h5052: y = 16'h200;
			16'h5053: y = 16'h200;
			16'h5054: y = 16'h200;
			16'h5055: y = 16'h200;
			16'h5056: y = 16'h200;
			16'h5057: y = 16'h200;
			16'h5058: y = 16'h200;
			16'h5059: y = 16'h200;
			16'h505a: y = 16'h200;
			16'h505b: y = 16'h200;
			16'h505c: y = 16'h200;
			16'h505d: y = 16'h200;
			16'h505e: y = 16'h200;
			16'h505f: y = 16'h200;
			16'h5060: y = 16'h200;
			16'h5061: y = 16'h200;
			16'h5062: y = 16'h200;
			16'h5063: y = 16'h200;
			16'h5064: y = 16'h200;
			16'h5065: y = 16'h200;
			16'h5066: y = 16'h200;
			16'h5067: y = 16'h200;
			16'h5068: y = 16'h200;
			16'h5069: y = 16'h200;
			16'h506a: y = 16'h200;
			16'h506b: y = 16'h200;
			16'h506c: y = 16'h200;
			16'h506d: y = 16'h200;
			16'h506e: y = 16'h200;
			16'h506f: y = 16'h200;
			16'h5070: y = 16'h200;
			16'h5071: y = 16'h200;
			16'h5072: y = 16'h200;
			16'h5073: y = 16'h200;
			16'h5074: y = 16'h200;
			16'h5075: y = 16'h200;
			16'h5076: y = 16'h200;
			16'h5077: y = 16'h200;
			16'h5078: y = 16'h200;
			16'h5079: y = 16'h200;
			16'h507a: y = 16'h200;
			16'h507b: y = 16'h200;
			16'h507c: y = 16'h200;
			16'h507d: y = 16'h200;
			16'h507e: y = 16'h200;
			16'h507f: y = 16'h200;
			16'h5080: y = 16'h200;
			16'h5081: y = 16'h200;
			16'h5082: y = 16'h200;
			16'h5083: y = 16'h200;
			16'h5084: y = 16'h200;
			16'h5085: y = 16'h200;
			16'h5086: y = 16'h200;
			16'h5087: y = 16'h200;
			16'h5088: y = 16'h200;
			16'h5089: y = 16'h200;
			16'h508a: y = 16'h200;
			16'h508b: y = 16'h200;
			16'h508c: y = 16'h200;
			16'h508d: y = 16'h200;
			16'h508e: y = 16'h200;
			16'h508f: y = 16'h200;
			16'h5090: y = 16'h200;
			16'h5091: y = 16'h200;
			16'h5092: y = 16'h200;
			16'h5093: y = 16'h200;
			16'h5094: y = 16'h200;
			16'h5095: y = 16'h200;
			16'h5096: y = 16'h200;
			16'h5097: y = 16'h200;
			16'h5098: y = 16'h200;
			16'h5099: y = 16'h200;
			16'h509a: y = 16'h200;
			16'h509b: y = 16'h200;
			16'h509c: y = 16'h200;
			16'h509d: y = 16'h200;
			16'h509e: y = 16'h200;
			16'h509f: y = 16'h200;
			16'h50a0: y = 16'h200;
			16'h50a1: y = 16'h200;
			16'h50a2: y = 16'h200;
			16'h50a3: y = 16'h200;
			16'h50a4: y = 16'h200;
			16'h50a5: y = 16'h200;
			16'h50a6: y = 16'h200;
			16'h50a7: y = 16'h200;
			16'h50a8: y = 16'h200;
			16'h50a9: y = 16'h200;
			16'h50aa: y = 16'h200;
			16'h50ab: y = 16'h200;
			16'h50ac: y = 16'h200;
			16'h50ad: y = 16'h200;
			16'h50ae: y = 16'h200;
			16'h50af: y = 16'h200;
			16'h50b0: y = 16'h200;
			16'h50b1: y = 16'h200;
			16'h50b2: y = 16'h200;
			16'h50b3: y = 16'h200;
			16'h50b4: y = 16'h200;
			16'h50b5: y = 16'h200;
			16'h50b6: y = 16'h200;
			16'h50b7: y = 16'h200;
			16'h50b8: y = 16'h200;
			16'h50b9: y = 16'h200;
			16'h50ba: y = 16'h200;
			16'h50bb: y = 16'h200;
			16'h50bc: y = 16'h200;
			16'h50bd: y = 16'h200;
			16'h50be: y = 16'h200;
			16'h50bf: y = 16'h200;
			16'h50c0: y = 16'h200;
			16'h50c1: y = 16'h200;
			16'h50c2: y = 16'h200;
			16'h50c3: y = 16'h200;
			16'h50c4: y = 16'h200;
			16'h50c5: y = 16'h200;
			16'h50c6: y = 16'h200;
			16'h50c7: y = 16'h200;
			16'h50c8: y = 16'h200;
			16'h50c9: y = 16'h200;
			16'h50ca: y = 16'h200;
			16'h50cb: y = 16'h200;
			16'h50cc: y = 16'h200;
			16'h50cd: y = 16'h200;
			16'h50ce: y = 16'h200;
			16'h50cf: y = 16'h200;
			16'h50d0: y = 16'h200;
			16'h50d1: y = 16'h200;
			16'h50d2: y = 16'h200;
			16'h50d3: y = 16'h200;
			16'h50d4: y = 16'h200;
			16'h50d5: y = 16'h200;
			16'h50d6: y = 16'h200;
			16'h50d7: y = 16'h200;
			16'h50d8: y = 16'h200;
			16'h50d9: y = 16'h200;
			16'h50da: y = 16'h200;
			16'h50db: y = 16'h200;
			16'h50dc: y = 16'h200;
			16'h50dd: y = 16'h200;
			16'h50de: y = 16'h200;
			16'h50df: y = 16'h200;
			16'h50e0: y = 16'h200;
			16'h50e1: y = 16'h200;
			16'h50e2: y = 16'h200;
			16'h50e3: y = 16'h200;
			16'h50e4: y = 16'h200;
			16'h50e5: y = 16'h200;
			16'h50e6: y = 16'h200;
			16'h50e7: y = 16'h200;
			16'h50e8: y = 16'h200;
			16'h50e9: y = 16'h200;
			16'h50ea: y = 16'h200;
			16'h50eb: y = 16'h200;
			16'h50ec: y = 16'h200;
			16'h50ed: y = 16'h200;
			16'h50ee: y = 16'h200;
			16'h50ef: y = 16'h200;
			16'h50f0: y = 16'h200;
			16'h50f1: y = 16'h200;
			16'h50f2: y = 16'h200;
			16'h50f3: y = 16'h200;
			16'h50f4: y = 16'h200;
			16'h50f5: y = 16'h200;
			16'h50f6: y = 16'h200;
			16'h50f7: y = 16'h200;
			16'h50f8: y = 16'h200;
			16'h50f9: y = 16'h200;
			16'h50fa: y = 16'h200;
			16'h50fb: y = 16'h200;
			16'h50fc: y = 16'h200;
			16'h50fd: y = 16'h200;
			16'h50fe: y = 16'h200;
			16'h50ff: y = 16'h200;
			16'h5100: y = 16'h200;
			16'h5101: y = 16'h200;
			16'h5102: y = 16'h200;
			16'h5103: y = 16'h200;
			16'h5104: y = 16'h200;
			16'h5105: y = 16'h200;
			16'h5106: y = 16'h200;
			16'h5107: y = 16'h200;
			16'h5108: y = 16'h200;
			16'h5109: y = 16'h200;
			16'h510a: y = 16'h200;
			16'h510b: y = 16'h200;
			16'h510c: y = 16'h200;
			16'h510d: y = 16'h200;
			16'h510e: y = 16'h200;
			16'h510f: y = 16'h200;
			16'h5110: y = 16'h200;
			16'h5111: y = 16'h200;
			16'h5112: y = 16'h200;
			16'h5113: y = 16'h200;
			16'h5114: y = 16'h200;
			16'h5115: y = 16'h200;
			16'h5116: y = 16'h200;
			16'h5117: y = 16'h200;
			16'h5118: y = 16'h200;
			16'h5119: y = 16'h200;
			16'h511a: y = 16'h200;
			16'h511b: y = 16'h200;
			16'h511c: y = 16'h200;
			16'h511d: y = 16'h200;
			16'h511e: y = 16'h200;
			16'h511f: y = 16'h200;
			16'h5120: y = 16'h200;
			16'h5121: y = 16'h200;
			16'h5122: y = 16'h200;
			16'h5123: y = 16'h200;
			16'h5124: y = 16'h200;
			16'h5125: y = 16'h200;
			16'h5126: y = 16'h200;
			16'h5127: y = 16'h200;
			16'h5128: y = 16'h200;
			16'h5129: y = 16'h200;
			16'h512a: y = 16'h200;
			16'h512b: y = 16'h200;
			16'h512c: y = 16'h200;
			16'h512d: y = 16'h200;
			16'h512e: y = 16'h200;
			16'h512f: y = 16'h200;
			16'h5130: y = 16'h200;
			16'h5131: y = 16'h200;
			16'h5132: y = 16'h200;
			16'h5133: y = 16'h200;
			16'h5134: y = 16'h200;
			16'h5135: y = 16'h200;
			16'h5136: y = 16'h200;
			16'h5137: y = 16'h200;
			16'h5138: y = 16'h200;
			16'h5139: y = 16'h200;
			16'h513a: y = 16'h200;
			16'h513b: y = 16'h200;
			16'h513c: y = 16'h200;
			16'h513d: y = 16'h200;
			16'h513e: y = 16'h200;
			16'h513f: y = 16'h200;
			16'h5140: y = 16'h200;
			16'h5141: y = 16'h200;
			16'h5142: y = 16'h200;
			16'h5143: y = 16'h200;
			16'h5144: y = 16'h200;
			16'h5145: y = 16'h200;
			16'h5146: y = 16'h200;
			16'h5147: y = 16'h200;
			16'h5148: y = 16'h200;
			16'h5149: y = 16'h200;
			16'h514a: y = 16'h200;
			16'h514b: y = 16'h200;
			16'h514c: y = 16'h200;
			16'h514d: y = 16'h200;
			16'h514e: y = 16'h200;
			16'h514f: y = 16'h200;
			16'h5150: y = 16'h200;
			16'h5151: y = 16'h200;
			16'h5152: y = 16'h200;
			16'h5153: y = 16'h200;
			16'h5154: y = 16'h200;
			16'h5155: y = 16'h200;
			16'h5156: y = 16'h200;
			16'h5157: y = 16'h200;
			16'h5158: y = 16'h200;
			16'h5159: y = 16'h200;
			16'h515a: y = 16'h200;
			16'h515b: y = 16'h200;
			16'h515c: y = 16'h200;
			16'h515d: y = 16'h200;
			16'h515e: y = 16'h200;
			16'h515f: y = 16'h200;
			16'h5160: y = 16'h200;
			16'h5161: y = 16'h200;
			16'h5162: y = 16'h200;
			16'h5163: y = 16'h200;
			16'h5164: y = 16'h200;
			16'h5165: y = 16'h200;
			16'h5166: y = 16'h200;
			16'h5167: y = 16'h200;
			16'h5168: y = 16'h200;
			16'h5169: y = 16'h200;
			16'h516a: y = 16'h200;
			16'h516b: y = 16'h200;
			16'h516c: y = 16'h200;
			16'h516d: y = 16'h200;
			16'h516e: y = 16'h200;
			16'h516f: y = 16'h200;
			16'h5170: y = 16'h200;
			16'h5171: y = 16'h200;
			16'h5172: y = 16'h200;
			16'h5173: y = 16'h200;
			16'h5174: y = 16'h200;
			16'h5175: y = 16'h200;
			16'h5176: y = 16'h200;
			16'h5177: y = 16'h200;
			16'h5178: y = 16'h200;
			16'h5179: y = 16'h200;
			16'h517a: y = 16'h200;
			16'h517b: y = 16'h200;
			16'h517c: y = 16'h200;
			16'h517d: y = 16'h200;
			16'h517e: y = 16'h200;
			16'h517f: y = 16'h200;
			16'h5180: y = 16'h200;
			16'h5181: y = 16'h200;
			16'h5182: y = 16'h200;
			16'h5183: y = 16'h200;
			16'h5184: y = 16'h200;
			16'h5185: y = 16'h200;
			16'h5186: y = 16'h200;
			16'h5187: y = 16'h200;
			16'h5188: y = 16'h200;
			16'h5189: y = 16'h200;
			16'h518a: y = 16'h200;
			16'h518b: y = 16'h200;
			16'h518c: y = 16'h200;
			16'h518d: y = 16'h200;
			16'h518e: y = 16'h200;
			16'h518f: y = 16'h200;
			16'h5190: y = 16'h200;
			16'h5191: y = 16'h200;
			16'h5192: y = 16'h200;
			16'h5193: y = 16'h200;
			16'h5194: y = 16'h200;
			16'h5195: y = 16'h200;
			16'h5196: y = 16'h200;
			16'h5197: y = 16'h200;
			16'h5198: y = 16'h200;
			16'h5199: y = 16'h200;
			16'h519a: y = 16'h200;
			16'h519b: y = 16'h200;
			16'h519c: y = 16'h200;
			16'h519d: y = 16'h200;
			16'h519e: y = 16'h200;
			16'h519f: y = 16'h200;
			16'h51a0: y = 16'h200;
			16'h51a1: y = 16'h200;
			16'h51a2: y = 16'h200;
			16'h51a3: y = 16'h200;
			16'h51a4: y = 16'h200;
			16'h51a5: y = 16'h200;
			16'h51a6: y = 16'h200;
			16'h51a7: y = 16'h200;
			16'h51a8: y = 16'h200;
			16'h51a9: y = 16'h200;
			16'h51aa: y = 16'h200;
			16'h51ab: y = 16'h200;
			16'h51ac: y = 16'h200;
			16'h51ad: y = 16'h200;
			16'h51ae: y = 16'h200;
			16'h51af: y = 16'h200;
			16'h51b0: y = 16'h200;
			16'h51b1: y = 16'h200;
			16'h51b2: y = 16'h200;
			16'h51b3: y = 16'h200;
			16'h51b4: y = 16'h200;
			16'h51b5: y = 16'h200;
			16'h51b6: y = 16'h200;
			16'h51b7: y = 16'h200;
			16'h51b8: y = 16'h200;
			16'h51b9: y = 16'h200;
			16'h51ba: y = 16'h200;
			16'h51bb: y = 16'h200;
			16'h51bc: y = 16'h200;
			16'h51bd: y = 16'h200;
			16'h51be: y = 16'h200;
			16'h51bf: y = 16'h200;
			16'h51c0: y = 16'h200;
			16'h51c1: y = 16'h200;
			16'h51c2: y = 16'h200;
			16'h51c3: y = 16'h200;
			16'h51c4: y = 16'h200;
			16'h51c5: y = 16'h200;
			16'h51c6: y = 16'h200;
			16'h51c7: y = 16'h200;
			16'h51c8: y = 16'h200;
			16'h51c9: y = 16'h200;
			16'h51ca: y = 16'h200;
			16'h51cb: y = 16'h200;
			16'h51cc: y = 16'h200;
			16'h51cd: y = 16'h200;
			16'h51ce: y = 16'h200;
			16'h51cf: y = 16'h200;
			16'h51d0: y = 16'h200;
			16'h51d1: y = 16'h200;
			16'h51d2: y = 16'h200;
			16'h51d3: y = 16'h200;
			16'h51d4: y = 16'h200;
			16'h51d5: y = 16'h200;
			16'h51d6: y = 16'h200;
			16'h51d7: y = 16'h200;
			16'h51d8: y = 16'h200;
			16'h51d9: y = 16'h200;
			16'h51da: y = 16'h200;
			16'h51db: y = 16'h200;
			16'h51dc: y = 16'h200;
			16'h51dd: y = 16'h200;
			16'h51de: y = 16'h200;
			16'h51df: y = 16'h200;
			16'h51e0: y = 16'h200;
			16'h51e1: y = 16'h200;
			16'h51e2: y = 16'h200;
			16'h51e3: y = 16'h200;
			16'h51e4: y = 16'h200;
			16'h51e5: y = 16'h200;
			16'h51e6: y = 16'h200;
			16'h51e7: y = 16'h200;
			16'h51e8: y = 16'h200;
			16'h51e9: y = 16'h200;
			16'h51ea: y = 16'h200;
			16'h51eb: y = 16'h200;
			16'h51ec: y = 16'h200;
			16'h51ed: y = 16'h200;
			16'h51ee: y = 16'h200;
			16'h51ef: y = 16'h200;
			16'h51f0: y = 16'h200;
			16'h51f1: y = 16'h200;
			16'h51f2: y = 16'h200;
			16'h51f3: y = 16'h200;
			16'h51f4: y = 16'h200;
			16'h51f5: y = 16'h200;
			16'h51f6: y = 16'h200;
			16'h51f7: y = 16'h200;
			16'h51f8: y = 16'h200;
			16'h51f9: y = 16'h200;
			16'h51fa: y = 16'h200;
			16'h51fb: y = 16'h200;
			16'h51fc: y = 16'h200;
			16'h51fd: y = 16'h200;
			16'h51fe: y = 16'h200;
			16'h51ff: y = 16'h200;
			16'h5200: y = 16'h200;
			16'h5201: y = 16'h200;
			16'h5202: y = 16'h200;
			16'h5203: y = 16'h200;
			16'h5204: y = 16'h200;
			16'h5205: y = 16'h200;
			16'h5206: y = 16'h200;
			16'h5207: y = 16'h200;
			16'h5208: y = 16'h200;
			16'h5209: y = 16'h200;
			16'h520a: y = 16'h200;
			16'h520b: y = 16'h200;
			16'h520c: y = 16'h200;
			16'h520d: y = 16'h200;
			16'h520e: y = 16'h200;
			16'h520f: y = 16'h200;
			16'h5210: y = 16'h200;
			16'h5211: y = 16'h200;
			16'h5212: y = 16'h200;
			16'h5213: y = 16'h200;
			16'h5214: y = 16'h200;
			16'h5215: y = 16'h200;
			16'h5216: y = 16'h200;
			16'h5217: y = 16'h200;
			16'h5218: y = 16'h200;
			16'h5219: y = 16'h200;
			16'h521a: y = 16'h200;
			16'h521b: y = 16'h200;
			16'h521c: y = 16'h200;
			16'h521d: y = 16'h200;
			16'h521e: y = 16'h200;
			16'h521f: y = 16'h200;
			16'h5220: y = 16'h200;
			16'h5221: y = 16'h200;
			16'h5222: y = 16'h200;
			16'h5223: y = 16'h200;
			16'h5224: y = 16'h200;
			16'h5225: y = 16'h200;
			16'h5226: y = 16'h200;
			16'h5227: y = 16'h200;
			16'h5228: y = 16'h200;
			16'h5229: y = 16'h200;
			16'h522a: y = 16'h200;
			16'h522b: y = 16'h200;
			16'h522c: y = 16'h200;
			16'h522d: y = 16'h200;
			16'h522e: y = 16'h200;
			16'h522f: y = 16'h200;
			16'h5230: y = 16'h200;
			16'h5231: y = 16'h200;
			16'h5232: y = 16'h200;
			16'h5233: y = 16'h200;
			16'h5234: y = 16'h200;
			16'h5235: y = 16'h200;
			16'h5236: y = 16'h200;
			16'h5237: y = 16'h200;
			16'h5238: y = 16'h200;
			16'h5239: y = 16'h200;
			16'h523a: y = 16'h200;
			16'h523b: y = 16'h200;
			16'h523c: y = 16'h200;
			16'h523d: y = 16'h200;
			16'h523e: y = 16'h200;
			16'h523f: y = 16'h200;
			16'h5240: y = 16'h200;
			16'h5241: y = 16'h200;
			16'h5242: y = 16'h200;
			16'h5243: y = 16'h200;
			16'h5244: y = 16'h200;
			16'h5245: y = 16'h200;
			16'h5246: y = 16'h200;
			16'h5247: y = 16'h200;
			16'h5248: y = 16'h200;
			16'h5249: y = 16'h200;
			16'h524a: y = 16'h200;
			16'h524b: y = 16'h200;
			16'h524c: y = 16'h200;
			16'h524d: y = 16'h200;
			16'h524e: y = 16'h200;
			16'h524f: y = 16'h200;
			16'h5250: y = 16'h200;
			16'h5251: y = 16'h200;
			16'h5252: y = 16'h200;
			16'h5253: y = 16'h200;
			16'h5254: y = 16'h200;
			16'h5255: y = 16'h200;
			16'h5256: y = 16'h200;
			16'h5257: y = 16'h200;
			16'h5258: y = 16'h200;
			16'h5259: y = 16'h200;
			16'h525a: y = 16'h200;
			16'h525b: y = 16'h200;
			16'h525c: y = 16'h200;
			16'h525d: y = 16'h200;
			16'h525e: y = 16'h200;
			16'h525f: y = 16'h200;
			16'h5260: y = 16'h200;
			16'h5261: y = 16'h200;
			16'h5262: y = 16'h200;
			16'h5263: y = 16'h200;
			16'h5264: y = 16'h200;
			16'h5265: y = 16'h200;
			16'h5266: y = 16'h200;
			16'h5267: y = 16'h200;
			16'h5268: y = 16'h200;
			16'h5269: y = 16'h200;
			16'h526a: y = 16'h200;
			16'h526b: y = 16'h200;
			16'h526c: y = 16'h200;
			16'h526d: y = 16'h200;
			16'h526e: y = 16'h200;
			16'h526f: y = 16'h200;
			16'h5270: y = 16'h200;
			16'h5271: y = 16'h200;
			16'h5272: y = 16'h200;
			16'h5273: y = 16'h200;
			16'h5274: y = 16'h200;
			16'h5275: y = 16'h200;
			16'h5276: y = 16'h200;
			16'h5277: y = 16'h200;
			16'h5278: y = 16'h200;
			16'h5279: y = 16'h200;
			16'h527a: y = 16'h200;
			16'h527b: y = 16'h200;
			16'h527c: y = 16'h200;
			16'h527d: y = 16'h200;
			16'h527e: y = 16'h200;
			16'h527f: y = 16'h200;
			16'h5280: y = 16'h200;
			16'h5281: y = 16'h200;
			16'h5282: y = 16'h200;
			16'h5283: y = 16'h200;
			16'h5284: y = 16'h200;
			16'h5285: y = 16'h200;
			16'h5286: y = 16'h200;
			16'h5287: y = 16'h200;
			16'h5288: y = 16'h200;
			16'h5289: y = 16'h200;
			16'h528a: y = 16'h200;
			16'h528b: y = 16'h200;
			16'h528c: y = 16'h200;
			16'h528d: y = 16'h200;
			16'h528e: y = 16'h200;
			16'h528f: y = 16'h200;
			16'h5290: y = 16'h200;
			16'h5291: y = 16'h200;
			16'h5292: y = 16'h200;
			16'h5293: y = 16'h200;
			16'h5294: y = 16'h200;
			16'h5295: y = 16'h200;
			16'h5296: y = 16'h200;
			16'h5297: y = 16'h200;
			16'h5298: y = 16'h200;
			16'h5299: y = 16'h200;
			16'h529a: y = 16'h200;
			16'h529b: y = 16'h200;
			16'h529c: y = 16'h200;
			16'h529d: y = 16'h200;
			16'h529e: y = 16'h200;
			16'h529f: y = 16'h200;
			16'h52a0: y = 16'h200;
			16'h52a1: y = 16'h200;
			16'h52a2: y = 16'h200;
			16'h52a3: y = 16'h200;
			16'h52a4: y = 16'h200;
			16'h52a5: y = 16'h200;
			16'h52a6: y = 16'h200;
			16'h52a7: y = 16'h200;
			16'h52a8: y = 16'h200;
			16'h52a9: y = 16'h200;
			16'h52aa: y = 16'h200;
			16'h52ab: y = 16'h200;
			16'h52ac: y = 16'h200;
			16'h52ad: y = 16'h200;
			16'h52ae: y = 16'h200;
			16'h52af: y = 16'h200;
			16'h52b0: y = 16'h200;
			16'h52b1: y = 16'h200;
			16'h52b2: y = 16'h200;
			16'h52b3: y = 16'h200;
			16'h52b4: y = 16'h200;
			16'h52b5: y = 16'h200;
			16'h52b6: y = 16'h200;
			16'h52b7: y = 16'h200;
			16'h52b8: y = 16'h200;
			16'h52b9: y = 16'h200;
			16'h52ba: y = 16'h200;
			16'h52bb: y = 16'h200;
			16'h52bc: y = 16'h200;
			16'h52bd: y = 16'h200;
			16'h52be: y = 16'h200;
			16'h52bf: y = 16'h200;
			16'h52c0: y = 16'h200;
			16'h52c1: y = 16'h200;
			16'h52c2: y = 16'h200;
			16'h52c3: y = 16'h200;
			16'h52c4: y = 16'h200;
			16'h52c5: y = 16'h200;
			16'h52c6: y = 16'h200;
			16'h52c7: y = 16'h200;
			16'h52c8: y = 16'h200;
			16'h52c9: y = 16'h200;
			16'h52ca: y = 16'h200;
			16'h52cb: y = 16'h200;
			16'h52cc: y = 16'h200;
			16'h52cd: y = 16'h200;
			16'h52ce: y = 16'h200;
			16'h52cf: y = 16'h200;
			16'h52d0: y = 16'h200;
			16'h52d1: y = 16'h200;
			16'h52d2: y = 16'h200;
			16'h52d3: y = 16'h200;
			16'h52d4: y = 16'h200;
			16'h52d5: y = 16'h200;
			16'h52d6: y = 16'h200;
			16'h52d7: y = 16'h200;
			16'h52d8: y = 16'h200;
			16'h52d9: y = 16'h200;
			16'h52da: y = 16'h200;
			16'h52db: y = 16'h200;
			16'h52dc: y = 16'h200;
			16'h52dd: y = 16'h200;
			16'h52de: y = 16'h200;
			16'h52df: y = 16'h200;
			16'h52e0: y = 16'h200;
			16'h52e1: y = 16'h200;
			16'h52e2: y = 16'h200;
			16'h52e3: y = 16'h200;
			16'h52e4: y = 16'h200;
			16'h52e5: y = 16'h200;
			16'h52e6: y = 16'h200;
			16'h52e7: y = 16'h200;
			16'h52e8: y = 16'h200;
			16'h52e9: y = 16'h200;
			16'h52ea: y = 16'h200;
			16'h52eb: y = 16'h200;
			16'h52ec: y = 16'h200;
			16'h52ed: y = 16'h200;
			16'h52ee: y = 16'h200;
			16'h52ef: y = 16'h200;
			16'h52f0: y = 16'h200;
			16'h52f1: y = 16'h200;
			16'h52f2: y = 16'h200;
			16'h52f3: y = 16'h200;
			16'h52f4: y = 16'h200;
			16'h52f5: y = 16'h200;
			16'h52f6: y = 16'h200;
			16'h52f7: y = 16'h200;
			16'h52f8: y = 16'h200;
			16'h52f9: y = 16'h200;
			16'h52fa: y = 16'h200;
			16'h52fb: y = 16'h200;
			16'h52fc: y = 16'h200;
			16'h52fd: y = 16'h200;
			16'h52fe: y = 16'h200;
			16'h52ff: y = 16'h200;
			16'h5300: y = 16'h200;
			16'h5301: y = 16'h200;
			16'h5302: y = 16'h200;
			16'h5303: y = 16'h200;
			16'h5304: y = 16'h200;
			16'h5305: y = 16'h200;
			16'h5306: y = 16'h200;
			16'h5307: y = 16'h200;
			16'h5308: y = 16'h200;
			16'h5309: y = 16'h200;
			16'h530a: y = 16'h200;
			16'h530b: y = 16'h200;
			16'h530c: y = 16'h200;
			16'h530d: y = 16'h200;
			16'h530e: y = 16'h200;
			16'h530f: y = 16'h200;
			16'h5310: y = 16'h200;
			16'h5311: y = 16'h200;
			16'h5312: y = 16'h200;
			16'h5313: y = 16'h200;
			16'h5314: y = 16'h200;
			16'h5315: y = 16'h200;
			16'h5316: y = 16'h200;
			16'h5317: y = 16'h200;
			16'h5318: y = 16'h200;
			16'h5319: y = 16'h200;
			16'h531a: y = 16'h200;
			16'h531b: y = 16'h200;
			16'h531c: y = 16'h200;
			16'h531d: y = 16'h200;
			16'h531e: y = 16'h200;
			16'h531f: y = 16'h200;
			16'h5320: y = 16'h200;
			16'h5321: y = 16'h200;
			16'h5322: y = 16'h200;
			16'h5323: y = 16'h200;
			16'h5324: y = 16'h200;
			16'h5325: y = 16'h200;
			16'h5326: y = 16'h200;
			16'h5327: y = 16'h200;
			16'h5328: y = 16'h200;
			16'h5329: y = 16'h200;
			16'h532a: y = 16'h200;
			16'h532b: y = 16'h200;
			16'h532c: y = 16'h200;
			16'h532d: y = 16'h200;
			16'h532e: y = 16'h200;
			16'h532f: y = 16'h200;
			16'h5330: y = 16'h200;
			16'h5331: y = 16'h200;
			16'h5332: y = 16'h200;
			16'h5333: y = 16'h200;
			16'h5334: y = 16'h200;
			16'h5335: y = 16'h200;
			16'h5336: y = 16'h200;
			16'h5337: y = 16'h200;
			16'h5338: y = 16'h200;
			16'h5339: y = 16'h200;
			16'h533a: y = 16'h200;
			16'h533b: y = 16'h200;
			16'h533c: y = 16'h200;
			16'h533d: y = 16'h200;
			16'h533e: y = 16'h200;
			16'h533f: y = 16'h200;
			16'h5340: y = 16'h200;
			16'h5341: y = 16'h200;
			16'h5342: y = 16'h200;
			16'h5343: y = 16'h200;
			16'h5344: y = 16'h200;
			16'h5345: y = 16'h200;
			16'h5346: y = 16'h200;
			16'h5347: y = 16'h200;
			16'h5348: y = 16'h200;
			16'h5349: y = 16'h200;
			16'h534a: y = 16'h200;
			16'h534b: y = 16'h200;
			16'h534c: y = 16'h200;
			16'h534d: y = 16'h200;
			16'h534e: y = 16'h200;
			16'h534f: y = 16'h200;
			16'h5350: y = 16'h200;
			16'h5351: y = 16'h200;
			16'h5352: y = 16'h200;
			16'h5353: y = 16'h200;
			16'h5354: y = 16'h200;
			16'h5355: y = 16'h200;
			16'h5356: y = 16'h200;
			16'h5357: y = 16'h200;
			16'h5358: y = 16'h200;
			16'h5359: y = 16'h200;
			16'h535a: y = 16'h200;
			16'h535b: y = 16'h200;
			16'h535c: y = 16'h200;
			16'h535d: y = 16'h200;
			16'h535e: y = 16'h200;
			16'h535f: y = 16'h200;
			16'h5360: y = 16'h200;
			16'h5361: y = 16'h200;
			16'h5362: y = 16'h200;
			16'h5363: y = 16'h200;
			16'h5364: y = 16'h200;
			16'h5365: y = 16'h200;
			16'h5366: y = 16'h200;
			16'h5367: y = 16'h200;
			16'h5368: y = 16'h200;
			16'h5369: y = 16'h200;
			16'h536a: y = 16'h200;
			16'h536b: y = 16'h200;
			16'h536c: y = 16'h200;
			16'h536d: y = 16'h200;
			16'h536e: y = 16'h200;
			16'h536f: y = 16'h200;
			16'h5370: y = 16'h200;
			16'h5371: y = 16'h200;
			16'h5372: y = 16'h200;
			16'h5373: y = 16'h200;
			16'h5374: y = 16'h200;
			16'h5375: y = 16'h200;
			16'h5376: y = 16'h200;
			16'h5377: y = 16'h200;
			16'h5378: y = 16'h200;
			16'h5379: y = 16'h200;
			16'h537a: y = 16'h200;
			16'h537b: y = 16'h200;
			16'h537c: y = 16'h200;
			16'h537d: y = 16'h200;
			16'h537e: y = 16'h200;
			16'h537f: y = 16'h200;
			16'h5380: y = 16'h200;
			16'h5381: y = 16'h200;
			16'h5382: y = 16'h200;
			16'h5383: y = 16'h200;
			16'h5384: y = 16'h200;
			16'h5385: y = 16'h200;
			16'h5386: y = 16'h200;
			16'h5387: y = 16'h200;
			16'h5388: y = 16'h200;
			16'h5389: y = 16'h200;
			16'h538a: y = 16'h200;
			16'h538b: y = 16'h200;
			16'h538c: y = 16'h200;
			16'h538d: y = 16'h200;
			16'h538e: y = 16'h200;
			16'h538f: y = 16'h200;
			16'h5390: y = 16'h200;
			16'h5391: y = 16'h200;
			16'h5392: y = 16'h200;
			16'h5393: y = 16'h200;
			16'h5394: y = 16'h200;
			16'h5395: y = 16'h200;
			16'h5396: y = 16'h200;
			16'h5397: y = 16'h200;
			16'h5398: y = 16'h200;
			16'h5399: y = 16'h200;
			16'h539a: y = 16'h200;
			16'h539b: y = 16'h200;
			16'h539c: y = 16'h200;
			16'h539d: y = 16'h200;
			16'h539e: y = 16'h200;
			16'h539f: y = 16'h200;
			16'h53a0: y = 16'h200;
			16'h53a1: y = 16'h200;
			16'h53a2: y = 16'h200;
			16'h53a3: y = 16'h200;
			16'h53a4: y = 16'h200;
			16'h53a5: y = 16'h200;
			16'h53a6: y = 16'h200;
			16'h53a7: y = 16'h200;
			16'h53a8: y = 16'h200;
			16'h53a9: y = 16'h200;
			16'h53aa: y = 16'h200;
			16'h53ab: y = 16'h200;
			16'h53ac: y = 16'h200;
			16'h53ad: y = 16'h200;
			16'h53ae: y = 16'h200;
			16'h53af: y = 16'h200;
			16'h53b0: y = 16'h200;
			16'h53b1: y = 16'h200;
			16'h53b2: y = 16'h200;
			16'h53b3: y = 16'h200;
			16'h53b4: y = 16'h200;
			16'h53b5: y = 16'h200;
			16'h53b6: y = 16'h200;
			16'h53b7: y = 16'h200;
			16'h53b8: y = 16'h200;
			16'h53b9: y = 16'h200;
			16'h53ba: y = 16'h200;
			16'h53bb: y = 16'h200;
			16'h53bc: y = 16'h200;
			16'h53bd: y = 16'h200;
			16'h53be: y = 16'h200;
			16'h53bf: y = 16'h200;
			16'h53c0: y = 16'h200;
			16'h53c1: y = 16'h200;
			16'h53c2: y = 16'h200;
			16'h53c3: y = 16'h200;
			16'h53c4: y = 16'h200;
			16'h53c5: y = 16'h200;
			16'h53c6: y = 16'h200;
			16'h53c7: y = 16'h200;
			16'h53c8: y = 16'h200;
			16'h53c9: y = 16'h200;
			16'h53ca: y = 16'h200;
			16'h53cb: y = 16'h200;
			16'h53cc: y = 16'h200;
			16'h53cd: y = 16'h200;
			16'h53ce: y = 16'h200;
			16'h53cf: y = 16'h200;
			16'h53d0: y = 16'h200;
			16'h53d1: y = 16'h200;
			16'h53d2: y = 16'h200;
			16'h53d3: y = 16'h200;
			16'h53d4: y = 16'h200;
			16'h53d5: y = 16'h200;
			16'h53d6: y = 16'h200;
			16'h53d7: y = 16'h200;
			16'h53d8: y = 16'h200;
			16'h53d9: y = 16'h200;
			16'h53da: y = 16'h200;
			16'h53db: y = 16'h200;
			16'h53dc: y = 16'h200;
			16'h53dd: y = 16'h200;
			16'h53de: y = 16'h200;
			16'h53df: y = 16'h200;
			16'h53e0: y = 16'h200;
			16'h53e1: y = 16'h200;
			16'h53e2: y = 16'h200;
			16'h53e3: y = 16'h200;
			16'h53e4: y = 16'h200;
			16'h53e5: y = 16'h200;
			16'h53e6: y = 16'h200;
			16'h53e7: y = 16'h200;
			16'h53e8: y = 16'h200;
			16'h53e9: y = 16'h200;
			16'h53ea: y = 16'h200;
			16'h53eb: y = 16'h200;
			16'h53ec: y = 16'h200;
			16'h53ed: y = 16'h200;
			16'h53ee: y = 16'h200;
			16'h53ef: y = 16'h200;
			16'h53f0: y = 16'h200;
			16'h53f1: y = 16'h200;
			16'h53f2: y = 16'h200;
			16'h53f3: y = 16'h200;
			16'h53f4: y = 16'h200;
			16'h53f5: y = 16'h200;
			16'h53f6: y = 16'h200;
			16'h53f7: y = 16'h200;
			16'h53f8: y = 16'h200;
			16'h53f9: y = 16'h200;
			16'h53fa: y = 16'h200;
			16'h53fb: y = 16'h200;
			16'h53fc: y = 16'h200;
			16'h53fd: y = 16'h200;
			16'h53fe: y = 16'h200;
			16'h53ff: y = 16'h200;
			16'h5400: y = 16'h200;
			16'h5401: y = 16'h200;
			16'h5402: y = 16'h200;
			16'h5403: y = 16'h200;
			16'h5404: y = 16'h200;
			16'h5405: y = 16'h200;
			16'h5406: y = 16'h200;
			16'h5407: y = 16'h200;
			16'h5408: y = 16'h200;
			16'h5409: y = 16'h200;
			16'h540a: y = 16'h200;
			16'h540b: y = 16'h200;
			16'h540c: y = 16'h200;
			16'h540d: y = 16'h200;
			16'h540e: y = 16'h200;
			16'h540f: y = 16'h200;
			16'h5410: y = 16'h200;
			16'h5411: y = 16'h200;
			16'h5412: y = 16'h200;
			16'h5413: y = 16'h200;
			16'h5414: y = 16'h200;
			16'h5415: y = 16'h200;
			16'h5416: y = 16'h200;
			16'h5417: y = 16'h200;
			16'h5418: y = 16'h200;
			16'h5419: y = 16'h200;
			16'h541a: y = 16'h200;
			16'h541b: y = 16'h200;
			16'h541c: y = 16'h200;
			16'h541d: y = 16'h200;
			16'h541e: y = 16'h200;
			16'h541f: y = 16'h200;
			16'h5420: y = 16'h200;
			16'h5421: y = 16'h200;
			16'h5422: y = 16'h200;
			16'h5423: y = 16'h200;
			16'h5424: y = 16'h200;
			16'h5425: y = 16'h200;
			16'h5426: y = 16'h200;
			16'h5427: y = 16'h200;
			16'h5428: y = 16'h200;
			16'h5429: y = 16'h200;
			16'h542a: y = 16'h200;
			16'h542b: y = 16'h200;
			16'h542c: y = 16'h200;
			16'h542d: y = 16'h200;
			16'h542e: y = 16'h200;
			16'h542f: y = 16'h200;
			16'h5430: y = 16'h200;
			16'h5431: y = 16'h200;
			16'h5432: y = 16'h200;
			16'h5433: y = 16'h200;
			16'h5434: y = 16'h200;
			16'h5435: y = 16'h200;
			16'h5436: y = 16'h200;
			16'h5437: y = 16'h200;
			16'h5438: y = 16'h200;
			16'h5439: y = 16'h200;
			16'h543a: y = 16'h200;
			16'h543b: y = 16'h200;
			16'h543c: y = 16'h200;
			16'h543d: y = 16'h200;
			16'h543e: y = 16'h200;
			16'h543f: y = 16'h200;
			16'h5440: y = 16'h200;
			16'h5441: y = 16'h200;
			16'h5442: y = 16'h200;
			16'h5443: y = 16'h200;
			16'h5444: y = 16'h200;
			16'h5445: y = 16'h200;
			16'h5446: y = 16'h200;
			16'h5447: y = 16'h200;
			16'h5448: y = 16'h200;
			16'h5449: y = 16'h200;
			16'h544a: y = 16'h200;
			16'h544b: y = 16'h200;
			16'h544c: y = 16'h200;
			16'h544d: y = 16'h200;
			16'h544e: y = 16'h200;
			16'h544f: y = 16'h200;
			16'h5450: y = 16'h200;
			16'h5451: y = 16'h200;
			16'h5452: y = 16'h200;
			16'h5453: y = 16'h200;
			16'h5454: y = 16'h200;
			16'h5455: y = 16'h200;
			16'h5456: y = 16'h200;
			16'h5457: y = 16'h200;
			16'h5458: y = 16'h200;
			16'h5459: y = 16'h200;
			16'h545a: y = 16'h200;
			16'h545b: y = 16'h200;
			16'h545c: y = 16'h200;
			16'h545d: y = 16'h200;
			16'h545e: y = 16'h200;
			16'h545f: y = 16'h200;
			16'h5460: y = 16'h200;
			16'h5461: y = 16'h200;
			16'h5462: y = 16'h200;
			16'h5463: y = 16'h200;
			16'h5464: y = 16'h200;
			16'h5465: y = 16'h200;
			16'h5466: y = 16'h200;
			16'h5467: y = 16'h200;
			16'h5468: y = 16'h200;
			16'h5469: y = 16'h200;
			16'h546a: y = 16'h200;
			16'h546b: y = 16'h200;
			16'h546c: y = 16'h200;
			16'h546d: y = 16'h200;
			16'h546e: y = 16'h200;
			16'h546f: y = 16'h200;
			16'h5470: y = 16'h200;
			16'h5471: y = 16'h200;
			16'h5472: y = 16'h200;
			16'h5473: y = 16'h200;
			16'h5474: y = 16'h200;
			16'h5475: y = 16'h200;
			16'h5476: y = 16'h200;
			16'h5477: y = 16'h200;
			16'h5478: y = 16'h200;
			16'h5479: y = 16'h200;
			16'h547a: y = 16'h200;
			16'h547b: y = 16'h200;
			16'h547c: y = 16'h200;
			16'h547d: y = 16'h200;
			16'h547e: y = 16'h200;
			16'h547f: y = 16'h200;
			16'h5480: y = 16'h200;
			16'h5481: y = 16'h200;
			16'h5482: y = 16'h200;
			16'h5483: y = 16'h200;
			16'h5484: y = 16'h200;
			16'h5485: y = 16'h200;
			16'h5486: y = 16'h200;
			16'h5487: y = 16'h200;
			16'h5488: y = 16'h200;
			16'h5489: y = 16'h200;
			16'h548a: y = 16'h200;
			16'h548b: y = 16'h200;
			16'h548c: y = 16'h200;
			16'h548d: y = 16'h200;
			16'h548e: y = 16'h200;
			16'h548f: y = 16'h200;
			16'h5490: y = 16'h200;
			16'h5491: y = 16'h200;
			16'h5492: y = 16'h200;
			16'h5493: y = 16'h200;
			16'h5494: y = 16'h200;
			16'h5495: y = 16'h200;
			16'h5496: y = 16'h200;
			16'h5497: y = 16'h200;
			16'h5498: y = 16'h200;
			16'h5499: y = 16'h200;
			16'h549a: y = 16'h200;
			16'h549b: y = 16'h200;
			16'h549c: y = 16'h200;
			16'h549d: y = 16'h200;
			16'h549e: y = 16'h200;
			16'h549f: y = 16'h200;
			16'h54a0: y = 16'h200;
			16'h54a1: y = 16'h200;
			16'h54a2: y = 16'h200;
			16'h54a3: y = 16'h200;
			16'h54a4: y = 16'h200;
			16'h54a5: y = 16'h200;
			16'h54a6: y = 16'h200;
			16'h54a7: y = 16'h200;
			16'h54a8: y = 16'h200;
			16'h54a9: y = 16'h200;
			16'h54aa: y = 16'h200;
			16'h54ab: y = 16'h200;
			16'h54ac: y = 16'h200;
			16'h54ad: y = 16'h200;
			16'h54ae: y = 16'h200;
			16'h54af: y = 16'h200;
			16'h54b0: y = 16'h200;
			16'h54b1: y = 16'h200;
			16'h54b2: y = 16'h200;
			16'h54b3: y = 16'h200;
			16'h54b4: y = 16'h200;
			16'h54b5: y = 16'h200;
			16'h54b6: y = 16'h200;
			16'h54b7: y = 16'h200;
			16'h54b8: y = 16'h200;
			16'h54b9: y = 16'h200;
			16'h54ba: y = 16'h200;
			16'h54bb: y = 16'h200;
			16'h54bc: y = 16'h200;
			16'h54bd: y = 16'h200;
			16'h54be: y = 16'h200;
			16'h54bf: y = 16'h200;
			16'h54c0: y = 16'h200;
			16'h54c1: y = 16'h200;
			16'h54c2: y = 16'h200;
			16'h54c3: y = 16'h200;
			16'h54c4: y = 16'h200;
			16'h54c5: y = 16'h200;
			16'h54c6: y = 16'h200;
			16'h54c7: y = 16'h200;
			16'h54c8: y = 16'h200;
			16'h54c9: y = 16'h200;
			16'h54ca: y = 16'h200;
			16'h54cb: y = 16'h200;
			16'h54cc: y = 16'h200;
			16'h54cd: y = 16'h200;
			16'h54ce: y = 16'h200;
			16'h54cf: y = 16'h200;
			16'h54d0: y = 16'h200;
			16'h54d1: y = 16'h200;
			16'h54d2: y = 16'h200;
			16'h54d3: y = 16'h200;
			16'h54d4: y = 16'h200;
			16'h54d5: y = 16'h200;
			16'h54d6: y = 16'h200;
			16'h54d7: y = 16'h200;
			16'h54d8: y = 16'h200;
			16'h54d9: y = 16'h200;
			16'h54da: y = 16'h200;
			16'h54db: y = 16'h200;
			16'h54dc: y = 16'h200;
			16'h54dd: y = 16'h200;
			16'h54de: y = 16'h200;
			16'h54df: y = 16'h200;
			16'h54e0: y = 16'h200;
			16'h54e1: y = 16'h200;
			16'h54e2: y = 16'h200;
			16'h54e3: y = 16'h200;
			16'h54e4: y = 16'h200;
			16'h54e5: y = 16'h200;
			16'h54e6: y = 16'h200;
			16'h54e7: y = 16'h200;
			16'h54e8: y = 16'h200;
			16'h54e9: y = 16'h200;
			16'h54ea: y = 16'h200;
			16'h54eb: y = 16'h200;
			16'h54ec: y = 16'h200;
			16'h54ed: y = 16'h200;
			16'h54ee: y = 16'h200;
			16'h54ef: y = 16'h200;
			16'h54f0: y = 16'h200;
			16'h54f1: y = 16'h200;
			16'h54f2: y = 16'h200;
			16'h54f3: y = 16'h200;
			16'h54f4: y = 16'h200;
			16'h54f5: y = 16'h200;
			16'h54f6: y = 16'h200;
			16'h54f7: y = 16'h200;
			16'h54f8: y = 16'h200;
			16'h54f9: y = 16'h200;
			16'h54fa: y = 16'h200;
			16'h54fb: y = 16'h200;
			16'h54fc: y = 16'h200;
			16'h54fd: y = 16'h200;
			16'h54fe: y = 16'h200;
			16'h54ff: y = 16'h200;
			16'h5500: y = 16'h200;
			16'h5501: y = 16'h200;
			16'h5502: y = 16'h200;
			16'h5503: y = 16'h200;
			16'h5504: y = 16'h200;
			16'h5505: y = 16'h200;
			16'h5506: y = 16'h200;
			16'h5507: y = 16'h200;
			16'h5508: y = 16'h200;
			16'h5509: y = 16'h200;
			16'h550a: y = 16'h200;
			16'h550b: y = 16'h200;
			16'h550c: y = 16'h200;
			16'h550d: y = 16'h200;
			16'h550e: y = 16'h200;
			16'h550f: y = 16'h200;
			16'h5510: y = 16'h200;
			16'h5511: y = 16'h200;
			16'h5512: y = 16'h200;
			16'h5513: y = 16'h200;
			16'h5514: y = 16'h200;
			16'h5515: y = 16'h200;
			16'h5516: y = 16'h200;
			16'h5517: y = 16'h200;
			16'h5518: y = 16'h200;
			16'h5519: y = 16'h200;
			16'h551a: y = 16'h200;
			16'h551b: y = 16'h200;
			16'h551c: y = 16'h200;
			16'h551d: y = 16'h200;
			16'h551e: y = 16'h200;
			16'h551f: y = 16'h200;
			16'h5520: y = 16'h200;
			16'h5521: y = 16'h200;
			16'h5522: y = 16'h200;
			16'h5523: y = 16'h200;
			16'h5524: y = 16'h200;
			16'h5525: y = 16'h200;
			16'h5526: y = 16'h200;
			16'h5527: y = 16'h200;
			16'h5528: y = 16'h200;
			16'h5529: y = 16'h200;
			16'h552a: y = 16'h200;
			16'h552b: y = 16'h200;
			16'h552c: y = 16'h200;
			16'h552d: y = 16'h200;
			16'h552e: y = 16'h200;
			16'h552f: y = 16'h200;
			16'h5530: y = 16'h200;
			16'h5531: y = 16'h200;
			16'h5532: y = 16'h200;
			16'h5533: y = 16'h200;
			16'h5534: y = 16'h200;
			16'h5535: y = 16'h200;
			16'h5536: y = 16'h200;
			16'h5537: y = 16'h200;
			16'h5538: y = 16'h200;
			16'h5539: y = 16'h200;
			16'h553a: y = 16'h200;
			16'h553b: y = 16'h200;
			16'h553c: y = 16'h200;
			16'h553d: y = 16'h200;
			16'h553e: y = 16'h200;
			16'h553f: y = 16'h200;
			16'h5540: y = 16'h200;
			16'h5541: y = 16'h200;
			16'h5542: y = 16'h200;
			16'h5543: y = 16'h200;
			16'h5544: y = 16'h200;
			16'h5545: y = 16'h200;
			16'h5546: y = 16'h200;
			16'h5547: y = 16'h200;
			16'h5548: y = 16'h200;
			16'h5549: y = 16'h200;
			16'h554a: y = 16'h200;
			16'h554b: y = 16'h200;
			16'h554c: y = 16'h200;
			16'h554d: y = 16'h200;
			16'h554e: y = 16'h200;
			16'h554f: y = 16'h200;
			16'h5550: y = 16'h200;
			16'h5551: y = 16'h200;
			16'h5552: y = 16'h200;
			16'h5553: y = 16'h200;
			16'h5554: y = 16'h200;
			16'h5555: y = 16'h200;
			16'h5556: y = 16'h200;
			16'h5557: y = 16'h200;
			16'h5558: y = 16'h200;
			16'h5559: y = 16'h200;
			16'h555a: y = 16'h200;
			16'h555b: y = 16'h200;
			16'h555c: y = 16'h200;
			16'h555d: y = 16'h200;
			16'h555e: y = 16'h200;
			16'h555f: y = 16'h200;
			16'h5560: y = 16'h200;
			16'h5561: y = 16'h200;
			16'h5562: y = 16'h200;
			16'h5563: y = 16'h200;
			16'h5564: y = 16'h200;
			16'h5565: y = 16'h200;
			16'h5566: y = 16'h200;
			16'h5567: y = 16'h200;
			16'h5568: y = 16'h200;
			16'h5569: y = 16'h200;
			16'h556a: y = 16'h200;
			16'h556b: y = 16'h200;
			16'h556c: y = 16'h200;
			16'h556d: y = 16'h200;
			16'h556e: y = 16'h200;
			16'h556f: y = 16'h200;
			16'h5570: y = 16'h200;
			16'h5571: y = 16'h200;
			16'h5572: y = 16'h200;
			16'h5573: y = 16'h200;
			16'h5574: y = 16'h200;
			16'h5575: y = 16'h200;
			16'h5576: y = 16'h200;
			16'h5577: y = 16'h200;
			16'h5578: y = 16'h200;
			16'h5579: y = 16'h200;
			16'h557a: y = 16'h200;
			16'h557b: y = 16'h200;
			16'h557c: y = 16'h200;
			16'h557d: y = 16'h200;
			16'h557e: y = 16'h200;
			16'h557f: y = 16'h200;
			16'h5580: y = 16'h200;
			16'h5581: y = 16'h200;
			16'h5582: y = 16'h200;
			16'h5583: y = 16'h200;
			16'h5584: y = 16'h200;
			16'h5585: y = 16'h200;
			16'h5586: y = 16'h200;
			16'h5587: y = 16'h200;
			16'h5588: y = 16'h200;
			16'h5589: y = 16'h200;
			16'h558a: y = 16'h200;
			16'h558b: y = 16'h200;
			16'h558c: y = 16'h200;
			16'h558d: y = 16'h200;
			16'h558e: y = 16'h200;
			16'h558f: y = 16'h200;
			16'h5590: y = 16'h200;
			16'h5591: y = 16'h200;
			16'h5592: y = 16'h200;
			16'h5593: y = 16'h200;
			16'h5594: y = 16'h200;
			16'h5595: y = 16'h200;
			16'h5596: y = 16'h200;
			16'h5597: y = 16'h200;
			16'h5598: y = 16'h200;
			16'h5599: y = 16'h200;
			16'h559a: y = 16'h200;
			16'h559b: y = 16'h200;
			16'h559c: y = 16'h200;
			16'h559d: y = 16'h200;
			16'h559e: y = 16'h200;
			16'h559f: y = 16'h200;
			16'h55a0: y = 16'h200;
			16'h55a1: y = 16'h200;
			16'h55a2: y = 16'h200;
			16'h55a3: y = 16'h200;
			16'h55a4: y = 16'h200;
			16'h55a5: y = 16'h200;
			16'h55a6: y = 16'h200;
			16'h55a7: y = 16'h200;
			16'h55a8: y = 16'h200;
			16'h55a9: y = 16'h200;
			16'h55aa: y = 16'h200;
			16'h55ab: y = 16'h200;
			16'h55ac: y = 16'h200;
			16'h55ad: y = 16'h200;
			16'h55ae: y = 16'h200;
			16'h55af: y = 16'h200;
			16'h55b0: y = 16'h200;
			16'h55b1: y = 16'h200;
			16'h55b2: y = 16'h200;
			16'h55b3: y = 16'h200;
			16'h55b4: y = 16'h200;
			16'h55b5: y = 16'h200;
			16'h55b6: y = 16'h200;
			16'h55b7: y = 16'h200;
			16'h55b8: y = 16'h200;
			16'h55b9: y = 16'h200;
			16'h55ba: y = 16'h200;
			16'h55bb: y = 16'h200;
			16'h55bc: y = 16'h200;
			16'h55bd: y = 16'h200;
			16'h55be: y = 16'h200;
			16'h55bf: y = 16'h200;
			16'h55c0: y = 16'h200;
			16'h55c1: y = 16'h200;
			16'h55c2: y = 16'h200;
			16'h55c3: y = 16'h200;
			16'h55c4: y = 16'h200;
			16'h55c5: y = 16'h200;
			16'h55c6: y = 16'h200;
			16'h55c7: y = 16'h200;
			16'h55c8: y = 16'h200;
			16'h55c9: y = 16'h200;
			16'h55ca: y = 16'h200;
			16'h55cb: y = 16'h200;
			16'h55cc: y = 16'h200;
			16'h55cd: y = 16'h200;
			16'h55ce: y = 16'h200;
			16'h55cf: y = 16'h200;
			16'h55d0: y = 16'h200;
			16'h55d1: y = 16'h200;
			16'h55d2: y = 16'h200;
			16'h55d3: y = 16'h200;
			16'h55d4: y = 16'h200;
			16'h55d5: y = 16'h200;
			16'h55d6: y = 16'h200;
			16'h55d7: y = 16'h200;
			16'h55d8: y = 16'h200;
			16'h55d9: y = 16'h200;
			16'h55da: y = 16'h200;
			16'h55db: y = 16'h200;
			16'h55dc: y = 16'h200;
			16'h55dd: y = 16'h200;
			16'h55de: y = 16'h200;
			16'h55df: y = 16'h200;
			16'h55e0: y = 16'h200;
			16'h55e1: y = 16'h200;
			16'h55e2: y = 16'h200;
			16'h55e3: y = 16'h200;
			16'h55e4: y = 16'h200;
			16'h55e5: y = 16'h200;
			16'h55e6: y = 16'h200;
			16'h55e7: y = 16'h200;
			16'h55e8: y = 16'h200;
			16'h55e9: y = 16'h200;
			16'h55ea: y = 16'h200;
			16'h55eb: y = 16'h200;
			16'h55ec: y = 16'h200;
			16'h55ed: y = 16'h200;
			16'h55ee: y = 16'h200;
			16'h55ef: y = 16'h200;
			16'h55f0: y = 16'h200;
			16'h55f1: y = 16'h200;
			16'h55f2: y = 16'h200;
			16'h55f3: y = 16'h200;
			16'h55f4: y = 16'h200;
			16'h55f5: y = 16'h200;
			16'h55f6: y = 16'h200;
			16'h55f7: y = 16'h200;
			16'h55f8: y = 16'h200;
			16'h55f9: y = 16'h200;
			16'h55fa: y = 16'h200;
			16'h55fb: y = 16'h200;
			16'h55fc: y = 16'h200;
			16'h55fd: y = 16'h200;
			16'h55fe: y = 16'h200;
			16'h55ff: y = 16'h200;
			16'h5600: y = 16'h200;
			16'h5601: y = 16'h200;
			16'h5602: y = 16'h200;
			16'h5603: y = 16'h200;
			16'h5604: y = 16'h200;
			16'h5605: y = 16'h200;
			16'h5606: y = 16'h200;
			16'h5607: y = 16'h200;
			16'h5608: y = 16'h200;
			16'h5609: y = 16'h200;
			16'h560a: y = 16'h200;
			16'h560b: y = 16'h200;
			16'h560c: y = 16'h200;
			16'h560d: y = 16'h200;
			16'h560e: y = 16'h200;
			16'h560f: y = 16'h200;
			16'h5610: y = 16'h200;
			16'h5611: y = 16'h200;
			16'h5612: y = 16'h200;
			16'h5613: y = 16'h200;
			16'h5614: y = 16'h200;
			16'h5615: y = 16'h200;
			16'h5616: y = 16'h200;
			16'h5617: y = 16'h200;
			16'h5618: y = 16'h200;
			16'h5619: y = 16'h200;
			16'h561a: y = 16'h200;
			16'h561b: y = 16'h200;
			16'h561c: y = 16'h200;
			16'h561d: y = 16'h200;
			16'h561e: y = 16'h200;
			16'h561f: y = 16'h200;
			16'h5620: y = 16'h200;
			16'h5621: y = 16'h200;
			16'h5622: y = 16'h200;
			16'h5623: y = 16'h200;
			16'h5624: y = 16'h200;
			16'h5625: y = 16'h200;
			16'h5626: y = 16'h200;
			16'h5627: y = 16'h200;
			16'h5628: y = 16'h200;
			16'h5629: y = 16'h200;
			16'h562a: y = 16'h200;
			16'h562b: y = 16'h200;
			16'h562c: y = 16'h200;
			16'h562d: y = 16'h200;
			16'h562e: y = 16'h200;
			16'h562f: y = 16'h200;
			16'h5630: y = 16'h200;
			16'h5631: y = 16'h200;
			16'h5632: y = 16'h200;
			16'h5633: y = 16'h200;
			16'h5634: y = 16'h200;
			16'h5635: y = 16'h200;
			16'h5636: y = 16'h200;
			16'h5637: y = 16'h200;
			16'h5638: y = 16'h200;
			16'h5639: y = 16'h200;
			16'h563a: y = 16'h200;
			16'h563b: y = 16'h200;
			16'h563c: y = 16'h200;
			16'h563d: y = 16'h200;
			16'h563e: y = 16'h200;
			16'h563f: y = 16'h200;
			16'h5640: y = 16'h200;
			16'h5641: y = 16'h200;
			16'h5642: y = 16'h200;
			16'h5643: y = 16'h200;
			16'h5644: y = 16'h200;
			16'h5645: y = 16'h200;
			16'h5646: y = 16'h200;
			16'h5647: y = 16'h200;
			16'h5648: y = 16'h200;
			16'h5649: y = 16'h200;
			16'h564a: y = 16'h200;
			16'h564b: y = 16'h200;
			16'h564c: y = 16'h200;
			16'h564d: y = 16'h200;
			16'h564e: y = 16'h200;
			16'h564f: y = 16'h200;
			16'h5650: y = 16'h200;
			16'h5651: y = 16'h200;
			16'h5652: y = 16'h200;
			16'h5653: y = 16'h200;
			16'h5654: y = 16'h200;
			16'h5655: y = 16'h200;
			16'h5656: y = 16'h200;
			16'h5657: y = 16'h200;
			16'h5658: y = 16'h200;
			16'h5659: y = 16'h200;
			16'h565a: y = 16'h200;
			16'h565b: y = 16'h200;
			16'h565c: y = 16'h200;
			16'h565d: y = 16'h200;
			16'h565e: y = 16'h200;
			16'h565f: y = 16'h200;
			16'h5660: y = 16'h200;
			16'h5661: y = 16'h200;
			16'h5662: y = 16'h200;
			16'h5663: y = 16'h200;
			16'h5664: y = 16'h200;
			16'h5665: y = 16'h200;
			16'h5666: y = 16'h200;
			16'h5667: y = 16'h200;
			16'h5668: y = 16'h200;
			16'h5669: y = 16'h200;
			16'h566a: y = 16'h200;
			16'h566b: y = 16'h200;
			16'h566c: y = 16'h200;
			16'h566d: y = 16'h200;
			16'h566e: y = 16'h200;
			16'h566f: y = 16'h200;
			16'h5670: y = 16'h200;
			16'h5671: y = 16'h200;
			16'h5672: y = 16'h200;
			16'h5673: y = 16'h200;
			16'h5674: y = 16'h200;
			16'h5675: y = 16'h200;
			16'h5676: y = 16'h200;
			16'h5677: y = 16'h200;
			16'h5678: y = 16'h200;
			16'h5679: y = 16'h200;
			16'h567a: y = 16'h200;
			16'h567b: y = 16'h200;
			16'h567c: y = 16'h200;
			16'h567d: y = 16'h200;
			16'h567e: y = 16'h200;
			16'h567f: y = 16'h200;
			16'h5680: y = 16'h200;
			16'h5681: y = 16'h200;
			16'h5682: y = 16'h200;
			16'h5683: y = 16'h200;
			16'h5684: y = 16'h200;
			16'h5685: y = 16'h200;
			16'h5686: y = 16'h200;
			16'h5687: y = 16'h200;
			16'h5688: y = 16'h200;
			16'h5689: y = 16'h200;
			16'h568a: y = 16'h200;
			16'h568b: y = 16'h200;
			16'h568c: y = 16'h200;
			16'h568d: y = 16'h200;
			16'h568e: y = 16'h200;
			16'h568f: y = 16'h200;
			16'h5690: y = 16'h200;
			16'h5691: y = 16'h200;
			16'h5692: y = 16'h200;
			16'h5693: y = 16'h200;
			16'h5694: y = 16'h200;
			16'h5695: y = 16'h200;
			16'h5696: y = 16'h200;
			16'h5697: y = 16'h200;
			16'h5698: y = 16'h200;
			16'h5699: y = 16'h200;
			16'h569a: y = 16'h200;
			16'h569b: y = 16'h200;
			16'h569c: y = 16'h200;
			16'h569d: y = 16'h200;
			16'h569e: y = 16'h200;
			16'h569f: y = 16'h200;
			16'h56a0: y = 16'h200;
			16'h56a1: y = 16'h200;
			16'h56a2: y = 16'h200;
			16'h56a3: y = 16'h200;
			16'h56a4: y = 16'h200;
			16'h56a5: y = 16'h200;
			16'h56a6: y = 16'h200;
			16'h56a7: y = 16'h200;
			16'h56a8: y = 16'h200;
			16'h56a9: y = 16'h200;
			16'h56aa: y = 16'h200;
			16'h56ab: y = 16'h200;
			16'h56ac: y = 16'h200;
			16'h56ad: y = 16'h200;
			16'h56ae: y = 16'h200;
			16'h56af: y = 16'h200;
			16'h56b0: y = 16'h200;
			16'h56b1: y = 16'h200;
			16'h56b2: y = 16'h200;
			16'h56b3: y = 16'h200;
			16'h56b4: y = 16'h200;
			16'h56b5: y = 16'h200;
			16'h56b6: y = 16'h200;
			16'h56b7: y = 16'h200;
			16'h56b8: y = 16'h200;
			16'h56b9: y = 16'h200;
			16'h56ba: y = 16'h200;
			16'h56bb: y = 16'h200;
			16'h56bc: y = 16'h200;
			16'h56bd: y = 16'h200;
			16'h56be: y = 16'h200;
			16'h56bf: y = 16'h200;
			16'h56c0: y = 16'h200;
			16'h56c1: y = 16'h200;
			16'h56c2: y = 16'h200;
			16'h56c3: y = 16'h200;
			16'h56c4: y = 16'h200;
			16'h56c5: y = 16'h200;
			16'h56c6: y = 16'h200;
			16'h56c7: y = 16'h200;
			16'h56c8: y = 16'h200;
			16'h56c9: y = 16'h200;
			16'h56ca: y = 16'h200;
			16'h56cb: y = 16'h200;
			16'h56cc: y = 16'h200;
			16'h56cd: y = 16'h200;
			16'h56ce: y = 16'h200;
			16'h56cf: y = 16'h200;
			16'h56d0: y = 16'h200;
			16'h56d1: y = 16'h200;
			16'h56d2: y = 16'h200;
			16'h56d3: y = 16'h200;
			16'h56d4: y = 16'h200;
			16'h56d5: y = 16'h200;
			16'h56d6: y = 16'h200;
			16'h56d7: y = 16'h200;
			16'h56d8: y = 16'h200;
			16'h56d9: y = 16'h200;
			16'h56da: y = 16'h200;
			16'h56db: y = 16'h200;
			16'h56dc: y = 16'h200;
			16'h56dd: y = 16'h200;
			16'h56de: y = 16'h200;
			16'h56df: y = 16'h200;
			16'h56e0: y = 16'h200;
			16'h56e1: y = 16'h200;
			16'h56e2: y = 16'h200;
			16'h56e3: y = 16'h200;
			16'h56e4: y = 16'h200;
			16'h56e5: y = 16'h200;
			16'h56e6: y = 16'h200;
			16'h56e7: y = 16'h200;
			16'h56e8: y = 16'h200;
			16'h56e9: y = 16'h200;
			16'h56ea: y = 16'h200;
			16'h56eb: y = 16'h200;
			16'h56ec: y = 16'h200;
			16'h56ed: y = 16'h200;
			16'h56ee: y = 16'h200;
			16'h56ef: y = 16'h200;
			16'h56f0: y = 16'h200;
			16'h56f1: y = 16'h200;
			16'h56f2: y = 16'h200;
			16'h56f3: y = 16'h200;
			16'h56f4: y = 16'h200;
			16'h56f5: y = 16'h200;
			16'h56f6: y = 16'h200;
			16'h56f7: y = 16'h200;
			16'h56f8: y = 16'h200;
			16'h56f9: y = 16'h200;
			16'h56fa: y = 16'h200;
			16'h56fb: y = 16'h200;
			16'h56fc: y = 16'h200;
			16'h56fd: y = 16'h200;
			16'h56fe: y = 16'h200;
			16'h56ff: y = 16'h200;
			16'h5700: y = 16'h200;
			16'h5701: y = 16'h200;
			16'h5702: y = 16'h200;
			16'h5703: y = 16'h200;
			16'h5704: y = 16'h200;
			16'h5705: y = 16'h200;
			16'h5706: y = 16'h200;
			16'h5707: y = 16'h200;
			16'h5708: y = 16'h200;
			16'h5709: y = 16'h200;
			16'h570a: y = 16'h200;
			16'h570b: y = 16'h200;
			16'h570c: y = 16'h200;
			16'h570d: y = 16'h200;
			16'h570e: y = 16'h200;
			16'h570f: y = 16'h200;
			16'h5710: y = 16'h200;
			16'h5711: y = 16'h200;
			16'h5712: y = 16'h200;
			16'h5713: y = 16'h200;
			16'h5714: y = 16'h200;
			16'h5715: y = 16'h200;
			16'h5716: y = 16'h200;
			16'h5717: y = 16'h200;
			16'h5718: y = 16'h200;
			16'h5719: y = 16'h200;
			16'h571a: y = 16'h200;
			16'h571b: y = 16'h200;
			16'h571c: y = 16'h200;
			16'h571d: y = 16'h200;
			16'h571e: y = 16'h200;
			16'h571f: y = 16'h200;
			16'h5720: y = 16'h200;
			16'h5721: y = 16'h200;
			16'h5722: y = 16'h200;
			16'h5723: y = 16'h200;
			16'h5724: y = 16'h200;
			16'h5725: y = 16'h200;
			16'h5726: y = 16'h200;
			16'h5727: y = 16'h200;
			16'h5728: y = 16'h200;
			16'h5729: y = 16'h200;
			16'h572a: y = 16'h200;
			16'h572b: y = 16'h200;
			16'h572c: y = 16'h200;
			16'h572d: y = 16'h200;
			16'h572e: y = 16'h200;
			16'h572f: y = 16'h200;
			16'h5730: y = 16'h200;
			16'h5731: y = 16'h200;
			16'h5732: y = 16'h200;
			16'h5733: y = 16'h200;
			16'h5734: y = 16'h200;
			16'h5735: y = 16'h200;
			16'h5736: y = 16'h200;
			16'h5737: y = 16'h200;
			16'h5738: y = 16'h200;
			16'h5739: y = 16'h200;
			16'h573a: y = 16'h200;
			16'h573b: y = 16'h200;
			16'h573c: y = 16'h200;
			16'h573d: y = 16'h200;
			16'h573e: y = 16'h200;
			16'h573f: y = 16'h200;
			16'h5740: y = 16'h200;
			16'h5741: y = 16'h200;
			16'h5742: y = 16'h200;
			16'h5743: y = 16'h200;
			16'h5744: y = 16'h200;
			16'h5745: y = 16'h200;
			16'h5746: y = 16'h200;
			16'h5747: y = 16'h200;
			16'h5748: y = 16'h200;
			16'h5749: y = 16'h200;
			16'h574a: y = 16'h200;
			16'h574b: y = 16'h200;
			16'h574c: y = 16'h200;
			16'h574d: y = 16'h200;
			16'h574e: y = 16'h200;
			16'h574f: y = 16'h200;
			16'h5750: y = 16'h200;
			16'h5751: y = 16'h200;
			16'h5752: y = 16'h200;
			16'h5753: y = 16'h200;
			16'h5754: y = 16'h200;
			16'h5755: y = 16'h200;
			16'h5756: y = 16'h200;
			16'h5757: y = 16'h200;
			16'h5758: y = 16'h200;
			16'h5759: y = 16'h200;
			16'h575a: y = 16'h200;
			16'h575b: y = 16'h200;
			16'h575c: y = 16'h200;
			16'h575d: y = 16'h200;
			16'h575e: y = 16'h200;
			16'h575f: y = 16'h200;
			16'h5760: y = 16'h200;
			16'h5761: y = 16'h200;
			16'h5762: y = 16'h200;
			16'h5763: y = 16'h200;
			16'h5764: y = 16'h200;
			16'h5765: y = 16'h200;
			16'h5766: y = 16'h200;
			16'h5767: y = 16'h200;
			16'h5768: y = 16'h200;
			16'h5769: y = 16'h200;
			16'h576a: y = 16'h200;
			16'h576b: y = 16'h200;
			16'h576c: y = 16'h200;
			16'h576d: y = 16'h200;
			16'h576e: y = 16'h200;
			16'h576f: y = 16'h200;
			16'h5770: y = 16'h200;
			16'h5771: y = 16'h200;
			16'h5772: y = 16'h200;
			16'h5773: y = 16'h200;
			16'h5774: y = 16'h200;
			16'h5775: y = 16'h200;
			16'h5776: y = 16'h200;
			16'h5777: y = 16'h200;
			16'h5778: y = 16'h200;
			16'h5779: y = 16'h200;
			16'h577a: y = 16'h200;
			16'h577b: y = 16'h200;
			16'h577c: y = 16'h200;
			16'h577d: y = 16'h200;
			16'h577e: y = 16'h200;
			16'h577f: y = 16'h200;
			16'h5780: y = 16'h200;
			16'h5781: y = 16'h200;
			16'h5782: y = 16'h200;
			16'h5783: y = 16'h200;
			16'h5784: y = 16'h200;
			16'h5785: y = 16'h200;
			16'h5786: y = 16'h200;
			16'h5787: y = 16'h200;
			16'h5788: y = 16'h200;
			16'h5789: y = 16'h200;
			16'h578a: y = 16'h200;
			16'h578b: y = 16'h200;
			16'h578c: y = 16'h200;
			16'h578d: y = 16'h200;
			16'h578e: y = 16'h200;
			16'h578f: y = 16'h200;
			16'h5790: y = 16'h200;
			16'h5791: y = 16'h200;
			16'h5792: y = 16'h200;
			16'h5793: y = 16'h200;
			16'h5794: y = 16'h200;
			16'h5795: y = 16'h200;
			16'h5796: y = 16'h200;
			16'h5797: y = 16'h200;
			16'h5798: y = 16'h200;
			16'h5799: y = 16'h200;
			16'h579a: y = 16'h200;
			16'h579b: y = 16'h200;
			16'h579c: y = 16'h200;
			16'h579d: y = 16'h200;
			16'h579e: y = 16'h200;
			16'h579f: y = 16'h200;
			16'h57a0: y = 16'h200;
			16'h57a1: y = 16'h200;
			16'h57a2: y = 16'h200;
			16'h57a3: y = 16'h200;
			16'h57a4: y = 16'h200;
			16'h57a5: y = 16'h200;
			16'h57a6: y = 16'h200;
			16'h57a7: y = 16'h200;
			16'h57a8: y = 16'h200;
			16'h57a9: y = 16'h200;
			16'h57aa: y = 16'h200;
			16'h57ab: y = 16'h200;
			16'h57ac: y = 16'h200;
			16'h57ad: y = 16'h200;
			16'h57ae: y = 16'h200;
			16'h57af: y = 16'h200;
			16'h57b0: y = 16'h200;
			16'h57b1: y = 16'h200;
			16'h57b2: y = 16'h200;
			16'h57b3: y = 16'h200;
			16'h57b4: y = 16'h200;
			16'h57b5: y = 16'h200;
			16'h57b6: y = 16'h200;
			16'h57b7: y = 16'h200;
			16'h57b8: y = 16'h200;
			16'h57b9: y = 16'h200;
			16'h57ba: y = 16'h200;
			16'h57bb: y = 16'h200;
			16'h57bc: y = 16'h200;
			16'h57bd: y = 16'h200;
			16'h57be: y = 16'h200;
			16'h57bf: y = 16'h200;
			16'h57c0: y = 16'h200;
			16'h57c1: y = 16'h200;
			16'h57c2: y = 16'h200;
			16'h57c3: y = 16'h200;
			16'h57c4: y = 16'h200;
			16'h57c5: y = 16'h200;
			16'h57c6: y = 16'h200;
			16'h57c7: y = 16'h200;
			16'h57c8: y = 16'h200;
			16'h57c9: y = 16'h200;
			16'h57ca: y = 16'h200;
			16'h57cb: y = 16'h200;
			16'h57cc: y = 16'h200;
			16'h57cd: y = 16'h200;
			16'h57ce: y = 16'h200;
			16'h57cf: y = 16'h200;
			16'h57d0: y = 16'h200;
			16'h57d1: y = 16'h200;
			16'h57d2: y = 16'h200;
			16'h57d3: y = 16'h200;
			16'h57d4: y = 16'h200;
			16'h57d5: y = 16'h200;
			16'h57d6: y = 16'h200;
			16'h57d7: y = 16'h200;
			16'h57d8: y = 16'h200;
			16'h57d9: y = 16'h200;
			16'h57da: y = 16'h200;
			16'h57db: y = 16'h200;
			16'h57dc: y = 16'h200;
			16'h57dd: y = 16'h200;
			16'h57de: y = 16'h200;
			16'h57df: y = 16'h200;
			16'h57e0: y = 16'h200;
			16'h57e1: y = 16'h200;
			16'h57e2: y = 16'h200;
			16'h57e3: y = 16'h200;
			16'h57e4: y = 16'h200;
			16'h57e5: y = 16'h200;
			16'h57e6: y = 16'h200;
			16'h57e7: y = 16'h200;
			16'h57e8: y = 16'h200;
			16'h57e9: y = 16'h200;
			16'h57ea: y = 16'h200;
			16'h57eb: y = 16'h200;
			16'h57ec: y = 16'h200;
			16'h57ed: y = 16'h200;
			16'h57ee: y = 16'h200;
			16'h57ef: y = 16'h200;
			16'h57f0: y = 16'h200;
			16'h57f1: y = 16'h200;
			16'h57f2: y = 16'h200;
			16'h57f3: y = 16'h200;
			16'h57f4: y = 16'h200;
			16'h57f5: y = 16'h200;
			16'h57f6: y = 16'h200;
			16'h57f7: y = 16'h200;
			16'h57f8: y = 16'h200;
			16'h57f9: y = 16'h200;
			16'h57fa: y = 16'h200;
			16'h57fb: y = 16'h200;
			16'h57fc: y = 16'h200;
			16'h57fd: y = 16'h200;
			16'h57fe: y = 16'h200;
			16'h57ff: y = 16'h200;
			16'h5800: y = 16'h200;
			16'h5801: y = 16'h200;
			16'h5802: y = 16'h200;
			16'h5803: y = 16'h200;
			16'h5804: y = 16'h200;
			16'h5805: y = 16'h200;
			16'h5806: y = 16'h200;
			16'h5807: y = 16'h200;
			16'h5808: y = 16'h200;
			16'h5809: y = 16'h200;
			16'h580a: y = 16'h200;
			16'h580b: y = 16'h200;
			16'h580c: y = 16'h200;
			16'h580d: y = 16'h200;
			16'h580e: y = 16'h200;
			16'h580f: y = 16'h200;
			16'h5810: y = 16'h200;
			16'h5811: y = 16'h200;
			16'h5812: y = 16'h200;
			16'h5813: y = 16'h200;
			16'h5814: y = 16'h200;
			16'h5815: y = 16'h200;
			16'h5816: y = 16'h200;
			16'h5817: y = 16'h200;
			16'h5818: y = 16'h200;
			16'h5819: y = 16'h200;
			16'h581a: y = 16'h200;
			16'h581b: y = 16'h200;
			16'h581c: y = 16'h200;
			16'h581d: y = 16'h200;
			16'h581e: y = 16'h200;
			16'h581f: y = 16'h200;
			16'h5820: y = 16'h200;
			16'h5821: y = 16'h200;
			16'h5822: y = 16'h200;
			16'h5823: y = 16'h200;
			16'h5824: y = 16'h200;
			16'h5825: y = 16'h200;
			16'h5826: y = 16'h200;
			16'h5827: y = 16'h200;
			16'h5828: y = 16'h200;
			16'h5829: y = 16'h200;
			16'h582a: y = 16'h200;
			16'h582b: y = 16'h200;
			16'h582c: y = 16'h200;
			16'h582d: y = 16'h200;
			16'h582e: y = 16'h200;
			16'h582f: y = 16'h200;
			16'h5830: y = 16'h200;
			16'h5831: y = 16'h200;
			16'h5832: y = 16'h200;
			16'h5833: y = 16'h200;
			16'h5834: y = 16'h200;
			16'h5835: y = 16'h200;
			16'h5836: y = 16'h200;
			16'h5837: y = 16'h200;
			16'h5838: y = 16'h200;
			16'h5839: y = 16'h200;
			16'h583a: y = 16'h200;
			16'h583b: y = 16'h200;
			16'h583c: y = 16'h200;
			16'h583d: y = 16'h200;
			16'h583e: y = 16'h200;
			16'h583f: y = 16'h200;
			16'h5840: y = 16'h200;
			16'h5841: y = 16'h200;
			16'h5842: y = 16'h200;
			16'h5843: y = 16'h200;
			16'h5844: y = 16'h200;
			16'h5845: y = 16'h200;
			16'h5846: y = 16'h200;
			16'h5847: y = 16'h200;
			16'h5848: y = 16'h200;
			16'h5849: y = 16'h200;
			16'h584a: y = 16'h200;
			16'h584b: y = 16'h200;
			16'h584c: y = 16'h200;
			16'h584d: y = 16'h200;
			16'h584e: y = 16'h200;
			16'h584f: y = 16'h200;
			16'h5850: y = 16'h200;
			16'h5851: y = 16'h200;
			16'h5852: y = 16'h200;
			16'h5853: y = 16'h200;
			16'h5854: y = 16'h200;
			16'h5855: y = 16'h200;
			16'h5856: y = 16'h200;
			16'h5857: y = 16'h200;
			16'h5858: y = 16'h200;
			16'h5859: y = 16'h200;
			16'h585a: y = 16'h200;
			16'h585b: y = 16'h200;
			16'h585c: y = 16'h200;
			16'h585d: y = 16'h200;
			16'h585e: y = 16'h200;
			16'h585f: y = 16'h200;
			16'h5860: y = 16'h200;
			16'h5861: y = 16'h200;
			16'h5862: y = 16'h200;
			16'h5863: y = 16'h200;
			16'h5864: y = 16'h200;
			16'h5865: y = 16'h200;
			16'h5866: y = 16'h200;
			16'h5867: y = 16'h200;
			16'h5868: y = 16'h200;
			16'h5869: y = 16'h200;
			16'h586a: y = 16'h200;
			16'h586b: y = 16'h200;
			16'h586c: y = 16'h200;
			16'h586d: y = 16'h200;
			16'h586e: y = 16'h200;
			16'h586f: y = 16'h200;
			16'h5870: y = 16'h200;
			16'h5871: y = 16'h200;
			16'h5872: y = 16'h200;
			16'h5873: y = 16'h200;
			16'h5874: y = 16'h200;
			16'h5875: y = 16'h200;
			16'h5876: y = 16'h200;
			16'h5877: y = 16'h200;
			16'h5878: y = 16'h200;
			16'h5879: y = 16'h200;
			16'h587a: y = 16'h200;
			16'h587b: y = 16'h200;
			16'h587c: y = 16'h200;
			16'h587d: y = 16'h200;
			16'h587e: y = 16'h200;
			16'h587f: y = 16'h200;
			16'h5880: y = 16'h200;
			16'h5881: y = 16'h200;
			16'h5882: y = 16'h200;
			16'h5883: y = 16'h200;
			16'h5884: y = 16'h200;
			16'h5885: y = 16'h200;
			16'h5886: y = 16'h200;
			16'h5887: y = 16'h200;
			16'h5888: y = 16'h200;
			16'h5889: y = 16'h200;
			16'h588a: y = 16'h200;
			16'h588b: y = 16'h200;
			16'h588c: y = 16'h200;
			16'h588d: y = 16'h200;
			16'h588e: y = 16'h200;
			16'h588f: y = 16'h200;
			16'h5890: y = 16'h200;
			16'h5891: y = 16'h200;
			16'h5892: y = 16'h200;
			16'h5893: y = 16'h200;
			16'h5894: y = 16'h200;
			16'h5895: y = 16'h200;
			16'h5896: y = 16'h200;
			16'h5897: y = 16'h200;
			16'h5898: y = 16'h200;
			16'h5899: y = 16'h200;
			16'h589a: y = 16'h200;
			16'h589b: y = 16'h200;
			16'h589c: y = 16'h200;
			16'h589d: y = 16'h200;
			16'h589e: y = 16'h200;
			16'h589f: y = 16'h200;
			16'h58a0: y = 16'h200;
			16'h58a1: y = 16'h200;
			16'h58a2: y = 16'h200;
			16'h58a3: y = 16'h200;
			16'h58a4: y = 16'h200;
			16'h58a5: y = 16'h200;
			16'h58a6: y = 16'h200;
			16'h58a7: y = 16'h200;
			16'h58a8: y = 16'h200;
			16'h58a9: y = 16'h200;
			16'h58aa: y = 16'h200;
			16'h58ab: y = 16'h200;
			16'h58ac: y = 16'h200;
			16'h58ad: y = 16'h200;
			16'h58ae: y = 16'h200;
			16'h58af: y = 16'h200;
			16'h58b0: y = 16'h200;
			16'h58b1: y = 16'h200;
			16'h58b2: y = 16'h200;
			16'h58b3: y = 16'h200;
			16'h58b4: y = 16'h200;
			16'h58b5: y = 16'h200;
			16'h58b6: y = 16'h200;
			16'h58b7: y = 16'h200;
			16'h58b8: y = 16'h200;
			16'h58b9: y = 16'h200;
			16'h58ba: y = 16'h200;
			16'h58bb: y = 16'h200;
			16'h58bc: y = 16'h200;
			16'h58bd: y = 16'h200;
			16'h58be: y = 16'h200;
			16'h58bf: y = 16'h200;
			16'h58c0: y = 16'h200;
			16'h58c1: y = 16'h200;
			16'h58c2: y = 16'h200;
			16'h58c3: y = 16'h200;
			16'h58c4: y = 16'h200;
			16'h58c5: y = 16'h200;
			16'h58c6: y = 16'h200;
			16'h58c7: y = 16'h200;
			16'h58c8: y = 16'h200;
			16'h58c9: y = 16'h200;
			16'h58ca: y = 16'h200;
			16'h58cb: y = 16'h200;
			16'h58cc: y = 16'h200;
			16'h58cd: y = 16'h200;
			16'h58ce: y = 16'h200;
			16'h58cf: y = 16'h200;
			16'h58d0: y = 16'h200;
			16'h58d1: y = 16'h200;
			16'h58d2: y = 16'h200;
			16'h58d3: y = 16'h200;
			16'h58d4: y = 16'h200;
			16'h58d5: y = 16'h200;
			16'h58d6: y = 16'h200;
			16'h58d7: y = 16'h200;
			16'h58d8: y = 16'h200;
			16'h58d9: y = 16'h200;
			16'h58da: y = 16'h200;
			16'h58db: y = 16'h200;
			16'h58dc: y = 16'h200;
			16'h58dd: y = 16'h200;
			16'h58de: y = 16'h200;
			16'h58df: y = 16'h200;
			16'h58e0: y = 16'h200;
			16'h58e1: y = 16'h200;
			16'h58e2: y = 16'h200;
			16'h58e3: y = 16'h200;
			16'h58e4: y = 16'h200;
			16'h58e5: y = 16'h200;
			16'h58e6: y = 16'h200;
			16'h58e7: y = 16'h200;
			16'h58e8: y = 16'h200;
			16'h58e9: y = 16'h200;
			16'h58ea: y = 16'h200;
			16'h58eb: y = 16'h200;
			16'h58ec: y = 16'h200;
			16'h58ed: y = 16'h200;
			16'h58ee: y = 16'h200;
			16'h58ef: y = 16'h200;
			16'h58f0: y = 16'h200;
			16'h58f1: y = 16'h200;
			16'h58f2: y = 16'h200;
			16'h58f3: y = 16'h200;
			16'h58f4: y = 16'h200;
			16'h58f5: y = 16'h200;
			16'h58f6: y = 16'h200;
			16'h58f7: y = 16'h200;
			16'h58f8: y = 16'h200;
			16'h58f9: y = 16'h200;
			16'h58fa: y = 16'h200;
			16'h58fb: y = 16'h200;
			16'h58fc: y = 16'h200;
			16'h58fd: y = 16'h200;
			16'h58fe: y = 16'h200;
			16'h58ff: y = 16'h200;
			16'h5900: y = 16'h200;
			16'h5901: y = 16'h200;
			16'h5902: y = 16'h200;
			16'h5903: y = 16'h200;
			16'h5904: y = 16'h200;
			16'h5905: y = 16'h200;
			16'h5906: y = 16'h200;
			16'h5907: y = 16'h200;
			16'h5908: y = 16'h200;
			16'h5909: y = 16'h200;
			16'h590a: y = 16'h200;
			16'h590b: y = 16'h200;
			16'h590c: y = 16'h200;
			16'h590d: y = 16'h200;
			16'h590e: y = 16'h200;
			16'h590f: y = 16'h200;
			16'h5910: y = 16'h200;
			16'h5911: y = 16'h200;
			16'h5912: y = 16'h200;
			16'h5913: y = 16'h200;
			16'h5914: y = 16'h200;
			16'h5915: y = 16'h200;
			16'h5916: y = 16'h200;
			16'h5917: y = 16'h200;
			16'h5918: y = 16'h200;
			16'h5919: y = 16'h200;
			16'h591a: y = 16'h200;
			16'h591b: y = 16'h200;
			16'h591c: y = 16'h200;
			16'h591d: y = 16'h200;
			16'h591e: y = 16'h200;
			16'h591f: y = 16'h200;
			16'h5920: y = 16'h200;
			16'h5921: y = 16'h200;
			16'h5922: y = 16'h200;
			16'h5923: y = 16'h200;
			16'h5924: y = 16'h200;
			16'h5925: y = 16'h200;
			16'h5926: y = 16'h200;
			16'h5927: y = 16'h200;
			16'h5928: y = 16'h200;
			16'h5929: y = 16'h200;
			16'h592a: y = 16'h200;
			16'h592b: y = 16'h200;
			16'h592c: y = 16'h200;
			16'h592d: y = 16'h200;
			16'h592e: y = 16'h200;
			16'h592f: y = 16'h200;
			16'h5930: y = 16'h200;
			16'h5931: y = 16'h200;
			16'h5932: y = 16'h200;
			16'h5933: y = 16'h200;
			16'h5934: y = 16'h200;
			16'h5935: y = 16'h200;
			16'h5936: y = 16'h200;
			16'h5937: y = 16'h200;
			16'h5938: y = 16'h200;
			16'h5939: y = 16'h200;
			16'h593a: y = 16'h200;
			16'h593b: y = 16'h200;
			16'h593c: y = 16'h200;
			16'h593d: y = 16'h200;
			16'h593e: y = 16'h200;
			16'h593f: y = 16'h200;
			16'h5940: y = 16'h200;
			16'h5941: y = 16'h200;
			16'h5942: y = 16'h200;
			16'h5943: y = 16'h200;
			16'h5944: y = 16'h200;
			16'h5945: y = 16'h200;
			16'h5946: y = 16'h200;
			16'h5947: y = 16'h200;
			16'h5948: y = 16'h200;
			16'h5949: y = 16'h200;
			16'h594a: y = 16'h200;
			16'h594b: y = 16'h200;
			16'h594c: y = 16'h200;
			16'h594d: y = 16'h200;
			16'h594e: y = 16'h200;
			16'h594f: y = 16'h200;
			16'h5950: y = 16'h200;
			16'h5951: y = 16'h200;
			16'h5952: y = 16'h200;
			16'h5953: y = 16'h200;
			16'h5954: y = 16'h200;
			16'h5955: y = 16'h200;
			16'h5956: y = 16'h200;
			16'h5957: y = 16'h200;
			16'h5958: y = 16'h200;
			16'h5959: y = 16'h200;
			16'h595a: y = 16'h200;
			16'h595b: y = 16'h200;
			16'h595c: y = 16'h200;
			16'h595d: y = 16'h200;
			16'h595e: y = 16'h200;
			16'h595f: y = 16'h200;
			16'h5960: y = 16'h200;
			16'h5961: y = 16'h200;
			16'h5962: y = 16'h200;
			16'h5963: y = 16'h200;
			16'h5964: y = 16'h200;
			16'h5965: y = 16'h200;
			16'h5966: y = 16'h200;
			16'h5967: y = 16'h200;
			16'h5968: y = 16'h200;
			16'h5969: y = 16'h200;
			16'h596a: y = 16'h200;
			16'h596b: y = 16'h200;
			16'h596c: y = 16'h200;
			16'h596d: y = 16'h200;
			16'h596e: y = 16'h200;
			16'h596f: y = 16'h200;
			16'h5970: y = 16'h200;
			16'h5971: y = 16'h200;
			16'h5972: y = 16'h200;
			16'h5973: y = 16'h200;
			16'h5974: y = 16'h200;
			16'h5975: y = 16'h200;
			16'h5976: y = 16'h200;
			16'h5977: y = 16'h200;
			16'h5978: y = 16'h200;
			16'h5979: y = 16'h200;
			16'h597a: y = 16'h200;
			16'h597b: y = 16'h200;
			16'h597c: y = 16'h200;
			16'h597d: y = 16'h200;
			16'h597e: y = 16'h200;
			16'h597f: y = 16'h200;
			16'h5980: y = 16'h200;
			16'h5981: y = 16'h200;
			16'h5982: y = 16'h200;
			16'h5983: y = 16'h200;
			16'h5984: y = 16'h200;
			16'h5985: y = 16'h200;
			16'h5986: y = 16'h200;
			16'h5987: y = 16'h200;
			16'h5988: y = 16'h200;
			16'h5989: y = 16'h200;
			16'h598a: y = 16'h200;
			16'h598b: y = 16'h200;
			16'h598c: y = 16'h200;
			16'h598d: y = 16'h200;
			16'h598e: y = 16'h200;
			16'h598f: y = 16'h200;
			16'h5990: y = 16'h200;
			16'h5991: y = 16'h200;
			16'h5992: y = 16'h200;
			16'h5993: y = 16'h200;
			16'h5994: y = 16'h200;
			16'h5995: y = 16'h200;
			16'h5996: y = 16'h200;
			16'h5997: y = 16'h200;
			16'h5998: y = 16'h200;
			16'h5999: y = 16'h200;
			16'h599a: y = 16'h200;
			16'h599b: y = 16'h200;
			16'h599c: y = 16'h200;
			16'h599d: y = 16'h200;
			16'h599e: y = 16'h200;
			16'h599f: y = 16'h200;
			16'h59a0: y = 16'h200;
			16'h59a1: y = 16'h200;
			16'h59a2: y = 16'h200;
			16'h59a3: y = 16'h200;
			16'h59a4: y = 16'h200;
			16'h59a5: y = 16'h200;
			16'h59a6: y = 16'h200;
			16'h59a7: y = 16'h200;
			16'h59a8: y = 16'h200;
			16'h59a9: y = 16'h200;
			16'h59aa: y = 16'h200;
			16'h59ab: y = 16'h200;
			16'h59ac: y = 16'h200;
			16'h59ad: y = 16'h200;
			16'h59ae: y = 16'h200;
			16'h59af: y = 16'h200;
			16'h59b0: y = 16'h200;
			16'h59b1: y = 16'h200;
			16'h59b2: y = 16'h200;
			16'h59b3: y = 16'h200;
			16'h59b4: y = 16'h200;
			16'h59b5: y = 16'h200;
			16'h59b6: y = 16'h200;
			16'h59b7: y = 16'h200;
			16'h59b8: y = 16'h200;
			16'h59b9: y = 16'h200;
			16'h59ba: y = 16'h200;
			16'h59bb: y = 16'h200;
			16'h59bc: y = 16'h200;
			16'h59bd: y = 16'h200;
			16'h59be: y = 16'h200;
			16'h59bf: y = 16'h200;
			16'h59c0: y = 16'h200;
			16'h59c1: y = 16'h200;
			16'h59c2: y = 16'h200;
			16'h59c3: y = 16'h200;
			16'h59c4: y = 16'h200;
			16'h59c5: y = 16'h200;
			16'h59c6: y = 16'h200;
			16'h59c7: y = 16'h200;
			16'h59c8: y = 16'h200;
			16'h59c9: y = 16'h200;
			16'h59ca: y = 16'h200;
			16'h59cb: y = 16'h200;
			16'h59cc: y = 16'h200;
			16'h59cd: y = 16'h200;
			16'h59ce: y = 16'h200;
			16'h59cf: y = 16'h200;
			16'h59d0: y = 16'h200;
			16'h59d1: y = 16'h200;
			16'h59d2: y = 16'h200;
			16'h59d3: y = 16'h200;
			16'h59d4: y = 16'h200;
			16'h59d5: y = 16'h200;
			16'h59d6: y = 16'h200;
			16'h59d7: y = 16'h200;
			16'h59d8: y = 16'h200;
			16'h59d9: y = 16'h200;
			16'h59da: y = 16'h200;
			16'h59db: y = 16'h200;
			16'h59dc: y = 16'h200;
			16'h59dd: y = 16'h200;
			16'h59de: y = 16'h200;
			16'h59df: y = 16'h200;
			16'h59e0: y = 16'h200;
			16'h59e1: y = 16'h200;
			16'h59e2: y = 16'h200;
			16'h59e3: y = 16'h200;
			16'h59e4: y = 16'h200;
			16'h59e5: y = 16'h200;
			16'h59e6: y = 16'h200;
			16'h59e7: y = 16'h200;
			16'h59e8: y = 16'h200;
			16'h59e9: y = 16'h200;
			16'h59ea: y = 16'h200;
			16'h59eb: y = 16'h200;
			16'h59ec: y = 16'h200;
			16'h59ed: y = 16'h200;
			16'h59ee: y = 16'h200;
			16'h59ef: y = 16'h200;
			16'h59f0: y = 16'h200;
			16'h59f1: y = 16'h200;
			16'h59f2: y = 16'h200;
			16'h59f3: y = 16'h200;
			16'h59f4: y = 16'h200;
			16'h59f5: y = 16'h200;
			16'h59f6: y = 16'h200;
			16'h59f7: y = 16'h200;
			16'h59f8: y = 16'h200;
			16'h59f9: y = 16'h200;
			16'h59fa: y = 16'h200;
			16'h59fb: y = 16'h200;
			16'h59fc: y = 16'h200;
			16'h59fd: y = 16'h200;
			16'h59fe: y = 16'h200;
			16'h59ff: y = 16'h200;
			16'h5a00: y = 16'h200;
			16'h5a01: y = 16'h200;
			16'h5a02: y = 16'h200;
			16'h5a03: y = 16'h200;
			16'h5a04: y = 16'h200;
			16'h5a05: y = 16'h200;
			16'h5a06: y = 16'h200;
			16'h5a07: y = 16'h200;
			16'h5a08: y = 16'h200;
			16'h5a09: y = 16'h200;
			16'h5a0a: y = 16'h200;
			16'h5a0b: y = 16'h200;
			16'h5a0c: y = 16'h200;
			16'h5a0d: y = 16'h200;
			16'h5a0e: y = 16'h200;
			16'h5a0f: y = 16'h200;
			16'h5a10: y = 16'h200;
			16'h5a11: y = 16'h200;
			16'h5a12: y = 16'h200;
			16'h5a13: y = 16'h200;
			16'h5a14: y = 16'h200;
			16'h5a15: y = 16'h200;
			16'h5a16: y = 16'h200;
			16'h5a17: y = 16'h200;
			16'h5a18: y = 16'h200;
			16'h5a19: y = 16'h200;
			16'h5a1a: y = 16'h200;
			16'h5a1b: y = 16'h200;
			16'h5a1c: y = 16'h200;
			16'h5a1d: y = 16'h200;
			16'h5a1e: y = 16'h200;
			16'h5a1f: y = 16'h200;
			16'h5a20: y = 16'h200;
			16'h5a21: y = 16'h200;
			16'h5a22: y = 16'h200;
			16'h5a23: y = 16'h200;
			16'h5a24: y = 16'h200;
			16'h5a25: y = 16'h200;
			16'h5a26: y = 16'h200;
			16'h5a27: y = 16'h200;
			16'h5a28: y = 16'h200;
			16'h5a29: y = 16'h200;
			16'h5a2a: y = 16'h200;
			16'h5a2b: y = 16'h200;
			16'h5a2c: y = 16'h200;
			16'h5a2d: y = 16'h200;
			16'h5a2e: y = 16'h200;
			16'h5a2f: y = 16'h200;
			16'h5a30: y = 16'h200;
			16'h5a31: y = 16'h200;
			16'h5a32: y = 16'h200;
			16'h5a33: y = 16'h200;
			16'h5a34: y = 16'h200;
			16'h5a35: y = 16'h200;
			16'h5a36: y = 16'h200;
			16'h5a37: y = 16'h200;
			16'h5a38: y = 16'h200;
			16'h5a39: y = 16'h200;
			16'h5a3a: y = 16'h200;
			16'h5a3b: y = 16'h200;
			16'h5a3c: y = 16'h200;
			16'h5a3d: y = 16'h200;
			16'h5a3e: y = 16'h200;
			16'h5a3f: y = 16'h200;
			16'h5a40: y = 16'h200;
			16'h5a41: y = 16'h200;
			16'h5a42: y = 16'h200;
			16'h5a43: y = 16'h200;
			16'h5a44: y = 16'h200;
			16'h5a45: y = 16'h200;
			16'h5a46: y = 16'h200;
			16'h5a47: y = 16'h200;
			16'h5a48: y = 16'h200;
			16'h5a49: y = 16'h200;
			16'h5a4a: y = 16'h200;
			16'h5a4b: y = 16'h200;
			16'h5a4c: y = 16'h200;
			16'h5a4d: y = 16'h200;
			16'h5a4e: y = 16'h200;
			16'h5a4f: y = 16'h200;
			16'h5a50: y = 16'h200;
			16'h5a51: y = 16'h200;
			16'h5a52: y = 16'h200;
			16'h5a53: y = 16'h200;
			16'h5a54: y = 16'h200;
			16'h5a55: y = 16'h200;
			16'h5a56: y = 16'h200;
			16'h5a57: y = 16'h200;
			16'h5a58: y = 16'h200;
			16'h5a59: y = 16'h200;
			16'h5a5a: y = 16'h200;
			16'h5a5b: y = 16'h200;
			16'h5a5c: y = 16'h200;
			16'h5a5d: y = 16'h200;
			16'h5a5e: y = 16'h200;
			16'h5a5f: y = 16'h200;
			16'h5a60: y = 16'h200;
			16'h5a61: y = 16'h200;
			16'h5a62: y = 16'h200;
			16'h5a63: y = 16'h200;
			16'h5a64: y = 16'h200;
			16'h5a65: y = 16'h200;
			16'h5a66: y = 16'h200;
			16'h5a67: y = 16'h200;
			16'h5a68: y = 16'h200;
			16'h5a69: y = 16'h200;
			16'h5a6a: y = 16'h200;
			16'h5a6b: y = 16'h200;
			16'h5a6c: y = 16'h200;
			16'h5a6d: y = 16'h200;
			16'h5a6e: y = 16'h200;
			16'h5a6f: y = 16'h200;
			16'h5a70: y = 16'h200;
			16'h5a71: y = 16'h200;
			16'h5a72: y = 16'h200;
			16'h5a73: y = 16'h200;
			16'h5a74: y = 16'h200;
			16'h5a75: y = 16'h200;
			16'h5a76: y = 16'h200;
			16'h5a77: y = 16'h200;
			16'h5a78: y = 16'h200;
			16'h5a79: y = 16'h200;
			16'h5a7a: y = 16'h200;
			16'h5a7b: y = 16'h200;
			16'h5a7c: y = 16'h200;
			16'h5a7d: y = 16'h200;
			16'h5a7e: y = 16'h200;
			16'h5a7f: y = 16'h200;
			16'h5a80: y = 16'h200;
			16'h5a81: y = 16'h200;
			16'h5a82: y = 16'h200;
			16'h5a83: y = 16'h200;
			16'h5a84: y = 16'h200;
			16'h5a85: y = 16'h200;
			16'h5a86: y = 16'h200;
			16'h5a87: y = 16'h200;
			16'h5a88: y = 16'h200;
			16'h5a89: y = 16'h200;
			16'h5a8a: y = 16'h200;
			16'h5a8b: y = 16'h200;
			16'h5a8c: y = 16'h200;
			16'h5a8d: y = 16'h200;
			16'h5a8e: y = 16'h200;
			16'h5a8f: y = 16'h200;
			16'h5a90: y = 16'h200;
			16'h5a91: y = 16'h200;
			16'h5a92: y = 16'h200;
			16'h5a93: y = 16'h200;
			16'h5a94: y = 16'h200;
			16'h5a95: y = 16'h200;
			16'h5a96: y = 16'h200;
			16'h5a97: y = 16'h200;
			16'h5a98: y = 16'h200;
			16'h5a99: y = 16'h200;
			16'h5a9a: y = 16'h200;
			16'h5a9b: y = 16'h200;
			16'h5a9c: y = 16'h200;
			16'h5a9d: y = 16'h200;
			16'h5a9e: y = 16'h200;
			16'h5a9f: y = 16'h200;
			16'h5aa0: y = 16'h200;
			16'h5aa1: y = 16'h200;
			16'h5aa2: y = 16'h200;
			16'h5aa3: y = 16'h200;
			16'h5aa4: y = 16'h200;
			16'h5aa5: y = 16'h200;
			16'h5aa6: y = 16'h200;
			16'h5aa7: y = 16'h200;
			16'h5aa8: y = 16'h200;
			16'h5aa9: y = 16'h200;
			16'h5aaa: y = 16'h200;
			16'h5aab: y = 16'h200;
			16'h5aac: y = 16'h200;
			16'h5aad: y = 16'h200;
			16'h5aae: y = 16'h200;
			16'h5aaf: y = 16'h200;
			16'h5ab0: y = 16'h200;
			16'h5ab1: y = 16'h200;
			16'h5ab2: y = 16'h200;
			16'h5ab3: y = 16'h200;
			16'h5ab4: y = 16'h200;
			16'h5ab5: y = 16'h200;
			16'h5ab6: y = 16'h200;
			16'h5ab7: y = 16'h200;
			16'h5ab8: y = 16'h200;
			16'h5ab9: y = 16'h200;
			16'h5aba: y = 16'h200;
			16'h5abb: y = 16'h200;
			16'h5abc: y = 16'h200;
			16'h5abd: y = 16'h200;
			16'h5abe: y = 16'h200;
			16'h5abf: y = 16'h200;
			16'h5ac0: y = 16'h200;
			16'h5ac1: y = 16'h200;
			16'h5ac2: y = 16'h200;
			16'h5ac3: y = 16'h200;
			16'h5ac4: y = 16'h200;
			16'h5ac5: y = 16'h200;
			16'h5ac6: y = 16'h200;
			16'h5ac7: y = 16'h200;
			16'h5ac8: y = 16'h200;
			16'h5ac9: y = 16'h200;
			16'h5aca: y = 16'h200;
			16'h5acb: y = 16'h200;
			16'h5acc: y = 16'h200;
			16'h5acd: y = 16'h200;
			16'h5ace: y = 16'h200;
			16'h5acf: y = 16'h200;
			16'h5ad0: y = 16'h200;
			16'h5ad1: y = 16'h200;
			16'h5ad2: y = 16'h200;
			16'h5ad3: y = 16'h200;
			16'h5ad4: y = 16'h200;
			16'h5ad5: y = 16'h200;
			16'h5ad6: y = 16'h200;
			16'h5ad7: y = 16'h200;
			16'h5ad8: y = 16'h200;
			16'h5ad9: y = 16'h200;
			16'h5ada: y = 16'h200;
			16'h5adb: y = 16'h200;
			16'h5adc: y = 16'h200;
			16'h5add: y = 16'h200;
			16'h5ade: y = 16'h200;
			16'h5adf: y = 16'h200;
			16'h5ae0: y = 16'h200;
			16'h5ae1: y = 16'h200;
			16'h5ae2: y = 16'h200;
			16'h5ae3: y = 16'h200;
			16'h5ae4: y = 16'h200;
			16'h5ae5: y = 16'h200;
			16'h5ae6: y = 16'h200;
			16'h5ae7: y = 16'h200;
			16'h5ae8: y = 16'h200;
			16'h5ae9: y = 16'h200;
			16'h5aea: y = 16'h200;
			16'h5aeb: y = 16'h200;
			16'h5aec: y = 16'h200;
			16'h5aed: y = 16'h200;
			16'h5aee: y = 16'h200;
			16'h5aef: y = 16'h200;
			16'h5af0: y = 16'h200;
			16'h5af1: y = 16'h200;
			16'h5af2: y = 16'h200;
			16'h5af3: y = 16'h200;
			16'h5af4: y = 16'h200;
			16'h5af5: y = 16'h200;
			16'h5af6: y = 16'h200;
			16'h5af7: y = 16'h200;
			16'h5af8: y = 16'h200;
			16'h5af9: y = 16'h200;
			16'h5afa: y = 16'h200;
			16'h5afb: y = 16'h200;
			16'h5afc: y = 16'h200;
			16'h5afd: y = 16'h200;
			16'h5afe: y = 16'h200;
			16'h5aff: y = 16'h200;
			16'h5b00: y = 16'h200;
			16'h5b01: y = 16'h200;
			16'h5b02: y = 16'h200;
			16'h5b03: y = 16'h200;
			16'h5b04: y = 16'h200;
			16'h5b05: y = 16'h200;
			16'h5b06: y = 16'h200;
			16'h5b07: y = 16'h200;
			16'h5b08: y = 16'h200;
			16'h5b09: y = 16'h200;
			16'h5b0a: y = 16'h200;
			16'h5b0b: y = 16'h200;
			16'h5b0c: y = 16'h200;
			16'h5b0d: y = 16'h200;
			16'h5b0e: y = 16'h200;
			16'h5b0f: y = 16'h200;
			16'h5b10: y = 16'h200;
			16'h5b11: y = 16'h200;
			16'h5b12: y = 16'h200;
			16'h5b13: y = 16'h200;
			16'h5b14: y = 16'h200;
			16'h5b15: y = 16'h200;
			16'h5b16: y = 16'h200;
			16'h5b17: y = 16'h200;
			16'h5b18: y = 16'h200;
			16'h5b19: y = 16'h200;
			16'h5b1a: y = 16'h200;
			16'h5b1b: y = 16'h200;
			16'h5b1c: y = 16'h200;
			16'h5b1d: y = 16'h200;
			16'h5b1e: y = 16'h200;
			16'h5b1f: y = 16'h200;
			16'h5b20: y = 16'h200;
			16'h5b21: y = 16'h200;
			16'h5b22: y = 16'h200;
			16'h5b23: y = 16'h200;
			16'h5b24: y = 16'h200;
			16'h5b25: y = 16'h200;
			16'h5b26: y = 16'h200;
			16'h5b27: y = 16'h200;
			16'h5b28: y = 16'h200;
			16'h5b29: y = 16'h200;
			16'h5b2a: y = 16'h200;
			16'h5b2b: y = 16'h200;
			16'h5b2c: y = 16'h200;
			16'h5b2d: y = 16'h200;
			16'h5b2e: y = 16'h200;
			16'h5b2f: y = 16'h200;
			16'h5b30: y = 16'h200;
			16'h5b31: y = 16'h200;
			16'h5b32: y = 16'h200;
			16'h5b33: y = 16'h200;
			16'h5b34: y = 16'h200;
			16'h5b35: y = 16'h200;
			16'h5b36: y = 16'h200;
			16'h5b37: y = 16'h200;
			16'h5b38: y = 16'h200;
			16'h5b39: y = 16'h200;
			16'h5b3a: y = 16'h200;
			16'h5b3b: y = 16'h200;
			16'h5b3c: y = 16'h200;
			16'h5b3d: y = 16'h200;
			16'h5b3e: y = 16'h200;
			16'h5b3f: y = 16'h200;
			16'h5b40: y = 16'h200;
			16'h5b41: y = 16'h200;
			16'h5b42: y = 16'h200;
			16'h5b43: y = 16'h200;
			16'h5b44: y = 16'h200;
			16'h5b45: y = 16'h200;
			16'h5b46: y = 16'h200;
			16'h5b47: y = 16'h200;
			16'h5b48: y = 16'h200;
			16'h5b49: y = 16'h200;
			16'h5b4a: y = 16'h200;
			16'h5b4b: y = 16'h200;
			16'h5b4c: y = 16'h200;
			16'h5b4d: y = 16'h200;
			16'h5b4e: y = 16'h200;
			16'h5b4f: y = 16'h200;
			16'h5b50: y = 16'h200;
			16'h5b51: y = 16'h200;
			16'h5b52: y = 16'h200;
			16'h5b53: y = 16'h200;
			16'h5b54: y = 16'h200;
			16'h5b55: y = 16'h200;
			16'h5b56: y = 16'h200;
			16'h5b57: y = 16'h200;
			16'h5b58: y = 16'h200;
			16'h5b59: y = 16'h200;
			16'h5b5a: y = 16'h200;
			16'h5b5b: y = 16'h200;
			16'h5b5c: y = 16'h200;
			16'h5b5d: y = 16'h200;
			16'h5b5e: y = 16'h200;
			16'h5b5f: y = 16'h200;
			16'h5b60: y = 16'h200;
			16'h5b61: y = 16'h200;
			16'h5b62: y = 16'h200;
			16'h5b63: y = 16'h200;
			16'h5b64: y = 16'h200;
			16'h5b65: y = 16'h200;
			16'h5b66: y = 16'h200;
			16'h5b67: y = 16'h200;
			16'h5b68: y = 16'h200;
			16'h5b69: y = 16'h200;
			16'h5b6a: y = 16'h200;
			16'h5b6b: y = 16'h200;
			16'h5b6c: y = 16'h200;
			16'h5b6d: y = 16'h200;
			16'h5b6e: y = 16'h200;
			16'h5b6f: y = 16'h200;
			16'h5b70: y = 16'h200;
			16'h5b71: y = 16'h200;
			16'h5b72: y = 16'h200;
			16'h5b73: y = 16'h200;
			16'h5b74: y = 16'h200;
			16'h5b75: y = 16'h200;
			16'h5b76: y = 16'h200;
			16'h5b77: y = 16'h200;
			16'h5b78: y = 16'h200;
			16'h5b79: y = 16'h200;
			16'h5b7a: y = 16'h200;
			16'h5b7b: y = 16'h200;
			16'h5b7c: y = 16'h200;
			16'h5b7d: y = 16'h200;
			16'h5b7e: y = 16'h200;
			16'h5b7f: y = 16'h200;
			16'h5b80: y = 16'h200;
			16'h5b81: y = 16'h200;
			16'h5b82: y = 16'h200;
			16'h5b83: y = 16'h200;
			16'h5b84: y = 16'h200;
			16'h5b85: y = 16'h200;
			16'h5b86: y = 16'h200;
			16'h5b87: y = 16'h200;
			16'h5b88: y = 16'h200;
			16'h5b89: y = 16'h200;
			16'h5b8a: y = 16'h200;
			16'h5b8b: y = 16'h200;
			16'h5b8c: y = 16'h200;
			16'h5b8d: y = 16'h200;
			16'h5b8e: y = 16'h200;
			16'h5b8f: y = 16'h200;
			16'h5b90: y = 16'h200;
			16'h5b91: y = 16'h200;
			16'h5b92: y = 16'h200;
			16'h5b93: y = 16'h200;
			16'h5b94: y = 16'h200;
			16'h5b95: y = 16'h200;
			16'h5b96: y = 16'h200;
			16'h5b97: y = 16'h200;
			16'h5b98: y = 16'h200;
			16'h5b99: y = 16'h200;
			16'h5b9a: y = 16'h200;
			16'h5b9b: y = 16'h200;
			16'h5b9c: y = 16'h200;
			16'h5b9d: y = 16'h200;
			16'h5b9e: y = 16'h200;
			16'h5b9f: y = 16'h200;
			16'h5ba0: y = 16'h200;
			16'h5ba1: y = 16'h200;
			16'h5ba2: y = 16'h200;
			16'h5ba3: y = 16'h200;
			16'h5ba4: y = 16'h200;
			16'h5ba5: y = 16'h200;
			16'h5ba6: y = 16'h200;
			16'h5ba7: y = 16'h200;
			16'h5ba8: y = 16'h200;
			16'h5ba9: y = 16'h200;
			16'h5baa: y = 16'h200;
			16'h5bab: y = 16'h200;
			16'h5bac: y = 16'h200;
			16'h5bad: y = 16'h200;
			16'h5bae: y = 16'h200;
			16'h5baf: y = 16'h200;
			16'h5bb0: y = 16'h200;
			16'h5bb1: y = 16'h200;
			16'h5bb2: y = 16'h200;
			16'h5bb3: y = 16'h200;
			16'h5bb4: y = 16'h200;
			16'h5bb5: y = 16'h200;
			16'h5bb6: y = 16'h200;
			16'h5bb7: y = 16'h200;
			16'h5bb8: y = 16'h200;
			16'h5bb9: y = 16'h200;
			16'h5bba: y = 16'h200;
			16'h5bbb: y = 16'h200;
			16'h5bbc: y = 16'h200;
			16'h5bbd: y = 16'h200;
			16'h5bbe: y = 16'h200;
			16'h5bbf: y = 16'h200;
			16'h5bc0: y = 16'h200;
			16'h5bc1: y = 16'h200;
			16'h5bc2: y = 16'h200;
			16'h5bc3: y = 16'h200;
			16'h5bc4: y = 16'h200;
			16'h5bc5: y = 16'h200;
			16'h5bc6: y = 16'h200;
			16'h5bc7: y = 16'h200;
			16'h5bc8: y = 16'h200;
			16'h5bc9: y = 16'h200;
			16'h5bca: y = 16'h200;
			16'h5bcb: y = 16'h200;
			16'h5bcc: y = 16'h200;
			16'h5bcd: y = 16'h200;
			16'h5bce: y = 16'h200;
			16'h5bcf: y = 16'h200;
			16'h5bd0: y = 16'h200;
			16'h5bd1: y = 16'h200;
			16'h5bd2: y = 16'h200;
			16'h5bd3: y = 16'h200;
			16'h5bd4: y = 16'h200;
			16'h5bd5: y = 16'h200;
			16'h5bd6: y = 16'h200;
			16'h5bd7: y = 16'h200;
			16'h5bd8: y = 16'h200;
			16'h5bd9: y = 16'h200;
			16'h5bda: y = 16'h200;
			16'h5bdb: y = 16'h200;
			16'h5bdc: y = 16'h200;
			16'h5bdd: y = 16'h200;
			16'h5bde: y = 16'h200;
			16'h5bdf: y = 16'h200;
			16'h5be0: y = 16'h200;
			16'h5be1: y = 16'h200;
			16'h5be2: y = 16'h200;
			16'h5be3: y = 16'h200;
			16'h5be4: y = 16'h200;
			16'h5be5: y = 16'h200;
			16'h5be6: y = 16'h200;
			16'h5be7: y = 16'h200;
			16'h5be8: y = 16'h200;
			16'h5be9: y = 16'h200;
			16'h5bea: y = 16'h200;
			16'h5beb: y = 16'h200;
			16'h5bec: y = 16'h200;
			16'h5bed: y = 16'h200;
			16'h5bee: y = 16'h200;
			16'h5bef: y = 16'h200;
			16'h5bf0: y = 16'h200;
			16'h5bf1: y = 16'h200;
			16'h5bf2: y = 16'h200;
			16'h5bf3: y = 16'h200;
			16'h5bf4: y = 16'h200;
			16'h5bf5: y = 16'h200;
			16'h5bf6: y = 16'h200;
			16'h5bf7: y = 16'h200;
			16'h5bf8: y = 16'h200;
			16'h5bf9: y = 16'h200;
			16'h5bfa: y = 16'h200;
			16'h5bfb: y = 16'h200;
			16'h5bfc: y = 16'h200;
			16'h5bfd: y = 16'h200;
			16'h5bfe: y = 16'h200;
			16'h5bff: y = 16'h200;
			16'h5c00: y = 16'h200;
			16'h5c01: y = 16'h200;
			16'h5c02: y = 16'h200;
			16'h5c03: y = 16'h200;
			16'h5c04: y = 16'h200;
			16'h5c05: y = 16'h200;
			16'h5c06: y = 16'h200;
			16'h5c07: y = 16'h200;
			16'h5c08: y = 16'h200;
			16'h5c09: y = 16'h200;
			16'h5c0a: y = 16'h200;
			16'h5c0b: y = 16'h200;
			16'h5c0c: y = 16'h200;
			16'h5c0d: y = 16'h200;
			16'h5c0e: y = 16'h200;
			16'h5c0f: y = 16'h200;
			16'h5c10: y = 16'h200;
			16'h5c11: y = 16'h200;
			16'h5c12: y = 16'h200;
			16'h5c13: y = 16'h200;
			16'h5c14: y = 16'h200;
			16'h5c15: y = 16'h200;
			16'h5c16: y = 16'h200;
			16'h5c17: y = 16'h200;
			16'h5c18: y = 16'h200;
			16'h5c19: y = 16'h200;
			16'h5c1a: y = 16'h200;
			16'h5c1b: y = 16'h200;
			16'h5c1c: y = 16'h200;
			16'h5c1d: y = 16'h200;
			16'h5c1e: y = 16'h200;
			16'h5c1f: y = 16'h200;
			16'h5c20: y = 16'h200;
			16'h5c21: y = 16'h200;
			16'h5c22: y = 16'h200;
			16'h5c23: y = 16'h200;
			16'h5c24: y = 16'h200;
			16'h5c25: y = 16'h200;
			16'h5c26: y = 16'h200;
			16'h5c27: y = 16'h200;
			16'h5c28: y = 16'h200;
			16'h5c29: y = 16'h200;
			16'h5c2a: y = 16'h200;
			16'h5c2b: y = 16'h200;
			16'h5c2c: y = 16'h200;
			16'h5c2d: y = 16'h200;
			16'h5c2e: y = 16'h200;
			16'h5c2f: y = 16'h200;
			16'h5c30: y = 16'h200;
			16'h5c31: y = 16'h200;
			16'h5c32: y = 16'h200;
			16'h5c33: y = 16'h200;
			16'h5c34: y = 16'h200;
			16'h5c35: y = 16'h200;
			16'h5c36: y = 16'h200;
			16'h5c37: y = 16'h200;
			16'h5c38: y = 16'h200;
			16'h5c39: y = 16'h200;
			16'h5c3a: y = 16'h200;
			16'h5c3b: y = 16'h200;
			16'h5c3c: y = 16'h200;
			16'h5c3d: y = 16'h200;
			16'h5c3e: y = 16'h200;
			16'h5c3f: y = 16'h200;
			16'h5c40: y = 16'h200;
			16'h5c41: y = 16'h200;
			16'h5c42: y = 16'h200;
			16'h5c43: y = 16'h200;
			16'h5c44: y = 16'h200;
			16'h5c45: y = 16'h200;
			16'h5c46: y = 16'h200;
			16'h5c47: y = 16'h200;
			16'h5c48: y = 16'h200;
			16'h5c49: y = 16'h200;
			16'h5c4a: y = 16'h200;
			16'h5c4b: y = 16'h200;
			16'h5c4c: y = 16'h200;
			16'h5c4d: y = 16'h200;
			16'h5c4e: y = 16'h200;
			16'h5c4f: y = 16'h200;
			16'h5c50: y = 16'h200;
			16'h5c51: y = 16'h200;
			16'h5c52: y = 16'h200;
			16'h5c53: y = 16'h200;
			16'h5c54: y = 16'h200;
			16'h5c55: y = 16'h200;
			16'h5c56: y = 16'h200;
			16'h5c57: y = 16'h200;
			16'h5c58: y = 16'h200;
			16'h5c59: y = 16'h200;
			16'h5c5a: y = 16'h200;
			16'h5c5b: y = 16'h200;
			16'h5c5c: y = 16'h200;
			16'h5c5d: y = 16'h200;
			16'h5c5e: y = 16'h200;
			16'h5c5f: y = 16'h200;
			16'h5c60: y = 16'h200;
			16'h5c61: y = 16'h200;
			16'h5c62: y = 16'h200;
			16'h5c63: y = 16'h200;
			16'h5c64: y = 16'h200;
			16'h5c65: y = 16'h200;
			16'h5c66: y = 16'h200;
			16'h5c67: y = 16'h200;
			16'h5c68: y = 16'h200;
			16'h5c69: y = 16'h200;
			16'h5c6a: y = 16'h200;
			16'h5c6b: y = 16'h200;
			16'h5c6c: y = 16'h200;
			16'h5c6d: y = 16'h200;
			16'h5c6e: y = 16'h200;
			16'h5c6f: y = 16'h200;
			16'h5c70: y = 16'h200;
			16'h5c71: y = 16'h200;
			16'h5c72: y = 16'h200;
			16'h5c73: y = 16'h200;
			16'h5c74: y = 16'h200;
			16'h5c75: y = 16'h200;
			16'h5c76: y = 16'h200;
			16'h5c77: y = 16'h200;
			16'h5c78: y = 16'h200;
			16'h5c79: y = 16'h200;
			16'h5c7a: y = 16'h200;
			16'h5c7b: y = 16'h200;
			16'h5c7c: y = 16'h200;
			16'h5c7d: y = 16'h200;
			16'h5c7e: y = 16'h200;
			16'h5c7f: y = 16'h200;
			16'h5c80: y = 16'h200;
			16'h5c81: y = 16'h200;
			16'h5c82: y = 16'h200;
			16'h5c83: y = 16'h200;
			16'h5c84: y = 16'h200;
			16'h5c85: y = 16'h200;
			16'h5c86: y = 16'h200;
			16'h5c87: y = 16'h200;
			16'h5c88: y = 16'h200;
			16'h5c89: y = 16'h200;
			16'h5c8a: y = 16'h200;
			16'h5c8b: y = 16'h200;
			16'h5c8c: y = 16'h200;
			16'h5c8d: y = 16'h200;
			16'h5c8e: y = 16'h200;
			16'h5c8f: y = 16'h200;
			16'h5c90: y = 16'h200;
			16'h5c91: y = 16'h200;
			16'h5c92: y = 16'h200;
			16'h5c93: y = 16'h200;
			16'h5c94: y = 16'h200;
			16'h5c95: y = 16'h200;
			16'h5c96: y = 16'h200;
			16'h5c97: y = 16'h200;
			16'h5c98: y = 16'h200;
			16'h5c99: y = 16'h200;
			16'h5c9a: y = 16'h200;
			16'h5c9b: y = 16'h200;
			16'h5c9c: y = 16'h200;
			16'h5c9d: y = 16'h200;
			16'h5c9e: y = 16'h200;
			16'h5c9f: y = 16'h200;
			16'h5ca0: y = 16'h200;
			16'h5ca1: y = 16'h200;
			16'h5ca2: y = 16'h200;
			16'h5ca3: y = 16'h200;
			16'h5ca4: y = 16'h200;
			16'h5ca5: y = 16'h200;
			16'h5ca6: y = 16'h200;
			16'h5ca7: y = 16'h200;
			16'h5ca8: y = 16'h200;
			16'h5ca9: y = 16'h200;
			16'h5caa: y = 16'h200;
			16'h5cab: y = 16'h200;
			16'h5cac: y = 16'h200;
			16'h5cad: y = 16'h200;
			16'h5cae: y = 16'h200;
			16'h5caf: y = 16'h200;
			16'h5cb0: y = 16'h200;
			16'h5cb1: y = 16'h200;
			16'h5cb2: y = 16'h200;
			16'h5cb3: y = 16'h200;
			16'h5cb4: y = 16'h200;
			16'h5cb5: y = 16'h200;
			16'h5cb6: y = 16'h200;
			16'h5cb7: y = 16'h200;
			16'h5cb8: y = 16'h200;
			16'h5cb9: y = 16'h200;
			16'h5cba: y = 16'h200;
			16'h5cbb: y = 16'h200;
			16'h5cbc: y = 16'h200;
			16'h5cbd: y = 16'h200;
			16'h5cbe: y = 16'h200;
			16'h5cbf: y = 16'h200;
			16'h5cc0: y = 16'h200;
			16'h5cc1: y = 16'h200;
			16'h5cc2: y = 16'h200;
			16'h5cc3: y = 16'h200;
			16'h5cc4: y = 16'h200;
			16'h5cc5: y = 16'h200;
			16'h5cc6: y = 16'h200;
			16'h5cc7: y = 16'h200;
			16'h5cc8: y = 16'h200;
			16'h5cc9: y = 16'h200;
			16'h5cca: y = 16'h200;
			16'h5ccb: y = 16'h200;
			16'h5ccc: y = 16'h200;
			16'h5ccd: y = 16'h200;
			16'h5cce: y = 16'h200;
			16'h5ccf: y = 16'h200;
			16'h5cd0: y = 16'h200;
			16'h5cd1: y = 16'h200;
			16'h5cd2: y = 16'h200;
			16'h5cd3: y = 16'h200;
			16'h5cd4: y = 16'h200;
			16'h5cd5: y = 16'h200;
			16'h5cd6: y = 16'h200;
			16'h5cd7: y = 16'h200;
			16'h5cd8: y = 16'h200;
			16'h5cd9: y = 16'h200;
			16'h5cda: y = 16'h200;
			16'h5cdb: y = 16'h200;
			16'h5cdc: y = 16'h200;
			16'h5cdd: y = 16'h200;
			16'h5cde: y = 16'h200;
			16'h5cdf: y = 16'h200;
			16'h5ce0: y = 16'h200;
			16'h5ce1: y = 16'h200;
			16'h5ce2: y = 16'h200;
			16'h5ce3: y = 16'h200;
			16'h5ce4: y = 16'h200;
			16'h5ce5: y = 16'h200;
			16'h5ce6: y = 16'h200;
			16'h5ce7: y = 16'h200;
			16'h5ce8: y = 16'h200;
			16'h5ce9: y = 16'h200;
			16'h5cea: y = 16'h200;
			16'h5ceb: y = 16'h200;
			16'h5cec: y = 16'h200;
			16'h5ced: y = 16'h200;
			16'h5cee: y = 16'h200;
			16'h5cef: y = 16'h200;
			16'h5cf0: y = 16'h200;
			16'h5cf1: y = 16'h200;
			16'h5cf2: y = 16'h200;
			16'h5cf3: y = 16'h200;
			16'h5cf4: y = 16'h200;
			16'h5cf5: y = 16'h200;
			16'h5cf6: y = 16'h200;
			16'h5cf7: y = 16'h200;
			16'h5cf8: y = 16'h200;
			16'h5cf9: y = 16'h200;
			16'h5cfa: y = 16'h200;
			16'h5cfb: y = 16'h200;
			16'h5cfc: y = 16'h200;
			16'h5cfd: y = 16'h200;
			16'h5cfe: y = 16'h200;
			16'h5cff: y = 16'h200;
			16'h5d00: y = 16'h200;
			16'h5d01: y = 16'h200;
			16'h5d02: y = 16'h200;
			16'h5d03: y = 16'h200;
			16'h5d04: y = 16'h200;
			16'h5d05: y = 16'h200;
			16'h5d06: y = 16'h200;
			16'h5d07: y = 16'h200;
			16'h5d08: y = 16'h200;
			16'h5d09: y = 16'h200;
			16'h5d0a: y = 16'h200;
			16'h5d0b: y = 16'h200;
			16'h5d0c: y = 16'h200;
			16'h5d0d: y = 16'h200;
			16'h5d0e: y = 16'h200;
			16'h5d0f: y = 16'h200;
			16'h5d10: y = 16'h200;
			16'h5d11: y = 16'h200;
			16'h5d12: y = 16'h200;
			16'h5d13: y = 16'h200;
			16'h5d14: y = 16'h200;
			16'h5d15: y = 16'h200;
			16'h5d16: y = 16'h200;
			16'h5d17: y = 16'h200;
			16'h5d18: y = 16'h200;
			16'h5d19: y = 16'h200;
			16'h5d1a: y = 16'h200;
			16'h5d1b: y = 16'h200;
			16'h5d1c: y = 16'h200;
			16'h5d1d: y = 16'h200;
			16'h5d1e: y = 16'h200;
			16'h5d1f: y = 16'h200;
			16'h5d20: y = 16'h200;
			16'h5d21: y = 16'h200;
			16'h5d22: y = 16'h200;
			16'h5d23: y = 16'h200;
			16'h5d24: y = 16'h200;
			16'h5d25: y = 16'h200;
			16'h5d26: y = 16'h200;
			16'h5d27: y = 16'h200;
			16'h5d28: y = 16'h200;
			16'h5d29: y = 16'h200;
			16'h5d2a: y = 16'h200;
			16'h5d2b: y = 16'h200;
			16'h5d2c: y = 16'h200;
			16'h5d2d: y = 16'h200;
			16'h5d2e: y = 16'h200;
			16'h5d2f: y = 16'h200;
			16'h5d30: y = 16'h200;
			16'h5d31: y = 16'h200;
			16'h5d32: y = 16'h200;
			16'h5d33: y = 16'h200;
			16'h5d34: y = 16'h200;
			16'h5d35: y = 16'h200;
			16'h5d36: y = 16'h200;
			16'h5d37: y = 16'h200;
			16'h5d38: y = 16'h200;
			16'h5d39: y = 16'h200;
			16'h5d3a: y = 16'h200;
			16'h5d3b: y = 16'h200;
			16'h5d3c: y = 16'h200;
			16'h5d3d: y = 16'h200;
			16'h5d3e: y = 16'h200;
			16'h5d3f: y = 16'h200;
			16'h5d40: y = 16'h200;
			16'h5d41: y = 16'h200;
			16'h5d42: y = 16'h200;
			16'h5d43: y = 16'h200;
			16'h5d44: y = 16'h200;
			16'h5d45: y = 16'h200;
			16'h5d46: y = 16'h200;
			16'h5d47: y = 16'h200;
			16'h5d48: y = 16'h200;
			16'h5d49: y = 16'h200;
			16'h5d4a: y = 16'h200;
			16'h5d4b: y = 16'h200;
			16'h5d4c: y = 16'h200;
			16'h5d4d: y = 16'h200;
			16'h5d4e: y = 16'h200;
			16'h5d4f: y = 16'h200;
			16'h5d50: y = 16'h200;
			16'h5d51: y = 16'h200;
			16'h5d52: y = 16'h200;
			16'h5d53: y = 16'h200;
			16'h5d54: y = 16'h200;
			16'h5d55: y = 16'h200;
			16'h5d56: y = 16'h200;
			16'h5d57: y = 16'h200;
			16'h5d58: y = 16'h200;
			16'h5d59: y = 16'h200;
			16'h5d5a: y = 16'h200;
			16'h5d5b: y = 16'h200;
			16'h5d5c: y = 16'h200;
			16'h5d5d: y = 16'h200;
			16'h5d5e: y = 16'h200;
			16'h5d5f: y = 16'h200;
			16'h5d60: y = 16'h200;
			16'h5d61: y = 16'h200;
			16'h5d62: y = 16'h200;
			16'h5d63: y = 16'h200;
			16'h5d64: y = 16'h200;
			16'h5d65: y = 16'h200;
			16'h5d66: y = 16'h200;
			16'h5d67: y = 16'h200;
			16'h5d68: y = 16'h200;
			16'h5d69: y = 16'h200;
			16'h5d6a: y = 16'h200;
			16'h5d6b: y = 16'h200;
			16'h5d6c: y = 16'h200;
			16'h5d6d: y = 16'h200;
			16'h5d6e: y = 16'h200;
			16'h5d6f: y = 16'h200;
			16'h5d70: y = 16'h200;
			16'h5d71: y = 16'h200;
			16'h5d72: y = 16'h200;
			16'h5d73: y = 16'h200;
			16'h5d74: y = 16'h200;
			16'h5d75: y = 16'h200;
			16'h5d76: y = 16'h200;
			16'h5d77: y = 16'h200;
			16'h5d78: y = 16'h200;
			16'h5d79: y = 16'h200;
			16'h5d7a: y = 16'h200;
			16'h5d7b: y = 16'h200;
			16'h5d7c: y = 16'h200;
			16'h5d7d: y = 16'h200;
			16'h5d7e: y = 16'h200;
			16'h5d7f: y = 16'h200;
			16'h5d80: y = 16'h200;
			16'h5d81: y = 16'h200;
			16'h5d82: y = 16'h200;
			16'h5d83: y = 16'h200;
			16'h5d84: y = 16'h200;
			16'h5d85: y = 16'h200;
			16'h5d86: y = 16'h200;
			16'h5d87: y = 16'h200;
			16'h5d88: y = 16'h200;
			16'h5d89: y = 16'h200;
			16'h5d8a: y = 16'h200;
			16'h5d8b: y = 16'h200;
			16'h5d8c: y = 16'h200;
			16'h5d8d: y = 16'h200;
			16'h5d8e: y = 16'h200;
			16'h5d8f: y = 16'h200;
			16'h5d90: y = 16'h200;
			16'h5d91: y = 16'h200;
			16'h5d92: y = 16'h200;
			16'h5d93: y = 16'h200;
			16'h5d94: y = 16'h200;
			16'h5d95: y = 16'h200;
			16'h5d96: y = 16'h200;
			16'h5d97: y = 16'h200;
			16'h5d98: y = 16'h200;
			16'h5d99: y = 16'h200;
			16'h5d9a: y = 16'h200;
			16'h5d9b: y = 16'h200;
			16'h5d9c: y = 16'h200;
			16'h5d9d: y = 16'h200;
			16'h5d9e: y = 16'h200;
			16'h5d9f: y = 16'h200;
			16'h5da0: y = 16'h200;
			16'h5da1: y = 16'h200;
			16'h5da2: y = 16'h200;
			16'h5da3: y = 16'h200;
			16'h5da4: y = 16'h200;
			16'h5da5: y = 16'h200;
			16'h5da6: y = 16'h200;
			16'h5da7: y = 16'h200;
			16'h5da8: y = 16'h200;
			16'h5da9: y = 16'h200;
			16'h5daa: y = 16'h200;
			16'h5dab: y = 16'h200;
			16'h5dac: y = 16'h200;
			16'h5dad: y = 16'h200;
			16'h5dae: y = 16'h200;
			16'h5daf: y = 16'h200;
			16'h5db0: y = 16'h200;
			16'h5db1: y = 16'h200;
			16'h5db2: y = 16'h200;
			16'h5db3: y = 16'h200;
			16'h5db4: y = 16'h200;
			16'h5db5: y = 16'h200;
			16'h5db6: y = 16'h200;
			16'h5db7: y = 16'h200;
			16'h5db8: y = 16'h200;
			16'h5db9: y = 16'h200;
			16'h5dba: y = 16'h200;
			16'h5dbb: y = 16'h200;
			16'h5dbc: y = 16'h200;
			16'h5dbd: y = 16'h200;
			16'h5dbe: y = 16'h200;
			16'h5dbf: y = 16'h200;
			16'h5dc0: y = 16'h200;
			16'h5dc1: y = 16'h200;
			16'h5dc2: y = 16'h200;
			16'h5dc3: y = 16'h200;
			16'h5dc4: y = 16'h200;
			16'h5dc5: y = 16'h200;
			16'h5dc6: y = 16'h200;
			16'h5dc7: y = 16'h200;
			16'h5dc8: y = 16'h200;
			16'h5dc9: y = 16'h200;
			16'h5dca: y = 16'h200;
			16'h5dcb: y = 16'h200;
			16'h5dcc: y = 16'h200;
			16'h5dcd: y = 16'h200;
			16'h5dce: y = 16'h200;
			16'h5dcf: y = 16'h200;
			16'h5dd0: y = 16'h200;
			16'h5dd1: y = 16'h200;
			16'h5dd2: y = 16'h200;
			16'h5dd3: y = 16'h200;
			16'h5dd4: y = 16'h200;
			16'h5dd5: y = 16'h200;
			16'h5dd6: y = 16'h200;
			16'h5dd7: y = 16'h200;
			16'h5dd8: y = 16'h200;
			16'h5dd9: y = 16'h200;
			16'h5dda: y = 16'h200;
			16'h5ddb: y = 16'h200;
			16'h5ddc: y = 16'h200;
			16'h5ddd: y = 16'h200;
			16'h5dde: y = 16'h200;
			16'h5ddf: y = 16'h200;
			16'h5de0: y = 16'h200;
			16'h5de1: y = 16'h200;
			16'h5de2: y = 16'h200;
			16'h5de3: y = 16'h200;
			16'h5de4: y = 16'h200;
			16'h5de5: y = 16'h200;
			16'h5de6: y = 16'h200;
			16'h5de7: y = 16'h200;
			16'h5de8: y = 16'h200;
			16'h5de9: y = 16'h200;
			16'h5dea: y = 16'h200;
			16'h5deb: y = 16'h200;
			16'h5dec: y = 16'h200;
			16'h5ded: y = 16'h200;
			16'h5dee: y = 16'h200;
			16'h5def: y = 16'h200;
			16'h5df0: y = 16'h200;
			16'h5df1: y = 16'h200;
			16'h5df2: y = 16'h200;
			16'h5df3: y = 16'h200;
			16'h5df4: y = 16'h200;
			16'h5df5: y = 16'h200;
			16'h5df6: y = 16'h200;
			16'h5df7: y = 16'h200;
			16'h5df8: y = 16'h200;
			16'h5df9: y = 16'h200;
			16'h5dfa: y = 16'h200;
			16'h5dfb: y = 16'h200;
			16'h5dfc: y = 16'h200;
			16'h5dfd: y = 16'h200;
			16'h5dfe: y = 16'h200;
			16'h5dff: y = 16'h200;
			16'h5e00: y = 16'h200;
			16'h5e01: y = 16'h200;
			16'h5e02: y = 16'h200;
			16'h5e03: y = 16'h200;
			16'h5e04: y = 16'h200;
			16'h5e05: y = 16'h200;
			16'h5e06: y = 16'h200;
			16'h5e07: y = 16'h200;
			16'h5e08: y = 16'h200;
			16'h5e09: y = 16'h200;
			16'h5e0a: y = 16'h200;
			16'h5e0b: y = 16'h200;
			16'h5e0c: y = 16'h200;
			16'h5e0d: y = 16'h200;
			16'h5e0e: y = 16'h200;
			16'h5e0f: y = 16'h200;
			16'h5e10: y = 16'h200;
			16'h5e11: y = 16'h200;
			16'h5e12: y = 16'h200;
			16'h5e13: y = 16'h200;
			16'h5e14: y = 16'h200;
			16'h5e15: y = 16'h200;
			16'h5e16: y = 16'h200;
			16'h5e17: y = 16'h200;
			16'h5e18: y = 16'h200;
			16'h5e19: y = 16'h200;
			16'h5e1a: y = 16'h200;
			16'h5e1b: y = 16'h200;
			16'h5e1c: y = 16'h200;
			16'h5e1d: y = 16'h200;
			16'h5e1e: y = 16'h200;
			16'h5e1f: y = 16'h200;
			16'h5e20: y = 16'h200;
			16'h5e21: y = 16'h200;
			16'h5e22: y = 16'h200;
			16'h5e23: y = 16'h200;
			16'h5e24: y = 16'h200;
			16'h5e25: y = 16'h200;
			16'h5e26: y = 16'h200;
			16'h5e27: y = 16'h200;
			16'h5e28: y = 16'h200;
			16'h5e29: y = 16'h200;
			16'h5e2a: y = 16'h200;
			16'h5e2b: y = 16'h200;
			16'h5e2c: y = 16'h200;
			16'h5e2d: y = 16'h200;
			16'h5e2e: y = 16'h200;
			16'h5e2f: y = 16'h200;
			16'h5e30: y = 16'h200;
			16'h5e31: y = 16'h200;
			16'h5e32: y = 16'h200;
			16'h5e33: y = 16'h200;
			16'h5e34: y = 16'h200;
			16'h5e35: y = 16'h200;
			16'h5e36: y = 16'h200;
			16'h5e37: y = 16'h200;
			16'h5e38: y = 16'h200;
			16'h5e39: y = 16'h200;
			16'h5e3a: y = 16'h200;
			16'h5e3b: y = 16'h200;
			16'h5e3c: y = 16'h200;
			16'h5e3d: y = 16'h200;
			16'h5e3e: y = 16'h200;
			16'h5e3f: y = 16'h200;
			16'h5e40: y = 16'h200;
			16'h5e41: y = 16'h200;
			16'h5e42: y = 16'h200;
			16'h5e43: y = 16'h200;
			16'h5e44: y = 16'h200;
			16'h5e45: y = 16'h200;
			16'h5e46: y = 16'h200;
			16'h5e47: y = 16'h200;
			16'h5e48: y = 16'h200;
			16'h5e49: y = 16'h200;
			16'h5e4a: y = 16'h200;
			16'h5e4b: y = 16'h200;
			16'h5e4c: y = 16'h200;
			16'h5e4d: y = 16'h200;
			16'h5e4e: y = 16'h200;
			16'h5e4f: y = 16'h200;
			16'h5e50: y = 16'h200;
			16'h5e51: y = 16'h200;
			16'h5e52: y = 16'h200;
			16'h5e53: y = 16'h200;
			16'h5e54: y = 16'h200;
			16'h5e55: y = 16'h200;
			16'h5e56: y = 16'h200;
			16'h5e57: y = 16'h200;
			16'h5e58: y = 16'h200;
			16'h5e59: y = 16'h200;
			16'h5e5a: y = 16'h200;
			16'h5e5b: y = 16'h200;
			16'h5e5c: y = 16'h200;
			16'h5e5d: y = 16'h200;
			16'h5e5e: y = 16'h200;
			16'h5e5f: y = 16'h200;
			16'h5e60: y = 16'h200;
			16'h5e61: y = 16'h200;
			16'h5e62: y = 16'h200;
			16'h5e63: y = 16'h200;
			16'h5e64: y = 16'h200;
			16'h5e65: y = 16'h200;
			16'h5e66: y = 16'h200;
			16'h5e67: y = 16'h200;
			16'h5e68: y = 16'h200;
			16'h5e69: y = 16'h200;
			16'h5e6a: y = 16'h200;
			16'h5e6b: y = 16'h200;
			16'h5e6c: y = 16'h200;
			16'h5e6d: y = 16'h200;
			16'h5e6e: y = 16'h200;
			16'h5e6f: y = 16'h200;
			16'h5e70: y = 16'h200;
			16'h5e71: y = 16'h200;
			16'h5e72: y = 16'h200;
			16'h5e73: y = 16'h200;
			16'h5e74: y = 16'h200;
			16'h5e75: y = 16'h200;
			16'h5e76: y = 16'h200;
			16'h5e77: y = 16'h200;
			16'h5e78: y = 16'h200;
			16'h5e79: y = 16'h200;
			16'h5e7a: y = 16'h200;
			16'h5e7b: y = 16'h200;
			16'h5e7c: y = 16'h200;
			16'h5e7d: y = 16'h200;
			16'h5e7e: y = 16'h200;
			16'h5e7f: y = 16'h200;
			16'h5e80: y = 16'h200;
			16'h5e81: y = 16'h200;
			16'h5e82: y = 16'h200;
			16'h5e83: y = 16'h200;
			16'h5e84: y = 16'h200;
			16'h5e85: y = 16'h200;
			16'h5e86: y = 16'h200;
			16'h5e87: y = 16'h200;
			16'h5e88: y = 16'h200;
			16'h5e89: y = 16'h200;
			16'h5e8a: y = 16'h200;
			16'h5e8b: y = 16'h200;
			16'h5e8c: y = 16'h200;
			16'h5e8d: y = 16'h200;
			16'h5e8e: y = 16'h200;
			16'h5e8f: y = 16'h200;
			16'h5e90: y = 16'h200;
			16'h5e91: y = 16'h200;
			16'h5e92: y = 16'h200;
			16'h5e93: y = 16'h200;
			16'h5e94: y = 16'h200;
			16'h5e95: y = 16'h200;
			16'h5e96: y = 16'h200;
			16'h5e97: y = 16'h200;
			16'h5e98: y = 16'h200;
			16'h5e99: y = 16'h200;
			16'h5e9a: y = 16'h200;
			16'h5e9b: y = 16'h200;
			16'h5e9c: y = 16'h200;
			16'h5e9d: y = 16'h200;
			16'h5e9e: y = 16'h200;
			16'h5e9f: y = 16'h200;
			16'h5ea0: y = 16'h200;
			16'h5ea1: y = 16'h200;
			16'h5ea2: y = 16'h200;
			16'h5ea3: y = 16'h200;
			16'h5ea4: y = 16'h200;
			16'h5ea5: y = 16'h200;
			16'h5ea6: y = 16'h200;
			16'h5ea7: y = 16'h200;
			16'h5ea8: y = 16'h200;
			16'h5ea9: y = 16'h200;
			16'h5eaa: y = 16'h200;
			16'h5eab: y = 16'h200;
			16'h5eac: y = 16'h200;
			16'h5ead: y = 16'h200;
			16'h5eae: y = 16'h200;
			16'h5eaf: y = 16'h200;
			16'h5eb0: y = 16'h200;
			16'h5eb1: y = 16'h200;
			16'h5eb2: y = 16'h200;
			16'h5eb3: y = 16'h200;
			16'h5eb4: y = 16'h200;
			16'h5eb5: y = 16'h200;
			16'h5eb6: y = 16'h200;
			16'h5eb7: y = 16'h200;
			16'h5eb8: y = 16'h200;
			16'h5eb9: y = 16'h200;
			16'h5eba: y = 16'h200;
			16'h5ebb: y = 16'h200;
			16'h5ebc: y = 16'h200;
			16'h5ebd: y = 16'h200;
			16'h5ebe: y = 16'h200;
			16'h5ebf: y = 16'h200;
			16'h5ec0: y = 16'h200;
			16'h5ec1: y = 16'h200;
			16'h5ec2: y = 16'h200;
			16'h5ec3: y = 16'h200;
			16'h5ec4: y = 16'h200;
			16'h5ec5: y = 16'h200;
			16'h5ec6: y = 16'h200;
			16'h5ec7: y = 16'h200;
			16'h5ec8: y = 16'h200;
			16'h5ec9: y = 16'h200;
			16'h5eca: y = 16'h200;
			16'h5ecb: y = 16'h200;
			16'h5ecc: y = 16'h200;
			16'h5ecd: y = 16'h200;
			16'h5ece: y = 16'h200;
			16'h5ecf: y = 16'h200;
			16'h5ed0: y = 16'h200;
			16'h5ed1: y = 16'h200;
			16'h5ed2: y = 16'h200;
			16'h5ed3: y = 16'h200;
			16'h5ed4: y = 16'h200;
			16'h5ed5: y = 16'h200;
			16'h5ed6: y = 16'h200;
			16'h5ed7: y = 16'h200;
			16'h5ed8: y = 16'h200;
			16'h5ed9: y = 16'h200;
			16'h5eda: y = 16'h200;
			16'h5edb: y = 16'h200;
			16'h5edc: y = 16'h200;
			16'h5edd: y = 16'h200;
			16'h5ede: y = 16'h200;
			16'h5edf: y = 16'h200;
			16'h5ee0: y = 16'h200;
			16'h5ee1: y = 16'h200;
			16'h5ee2: y = 16'h200;
			16'h5ee3: y = 16'h200;
			16'h5ee4: y = 16'h200;
			16'h5ee5: y = 16'h200;
			16'h5ee6: y = 16'h200;
			16'h5ee7: y = 16'h200;
			16'h5ee8: y = 16'h200;
			16'h5ee9: y = 16'h200;
			16'h5eea: y = 16'h200;
			16'h5eeb: y = 16'h200;
			16'h5eec: y = 16'h200;
			16'h5eed: y = 16'h200;
			16'h5eee: y = 16'h200;
			16'h5eef: y = 16'h200;
			16'h5ef0: y = 16'h200;
			16'h5ef1: y = 16'h200;
			16'h5ef2: y = 16'h200;
			16'h5ef3: y = 16'h200;
			16'h5ef4: y = 16'h200;
			16'h5ef5: y = 16'h200;
			16'h5ef6: y = 16'h200;
			16'h5ef7: y = 16'h200;
			16'h5ef8: y = 16'h200;
			16'h5ef9: y = 16'h200;
			16'h5efa: y = 16'h200;
			16'h5efb: y = 16'h200;
			16'h5efc: y = 16'h200;
			16'h5efd: y = 16'h200;
			16'h5efe: y = 16'h200;
			16'h5eff: y = 16'h200;
			16'h5f00: y = 16'h200;
			16'h5f01: y = 16'h200;
			16'h5f02: y = 16'h200;
			16'h5f03: y = 16'h200;
			16'h5f04: y = 16'h200;
			16'h5f05: y = 16'h200;
			16'h5f06: y = 16'h200;
			16'h5f07: y = 16'h200;
			16'h5f08: y = 16'h200;
			16'h5f09: y = 16'h200;
			16'h5f0a: y = 16'h200;
			16'h5f0b: y = 16'h200;
			16'h5f0c: y = 16'h200;
			16'h5f0d: y = 16'h200;
			16'h5f0e: y = 16'h200;
			16'h5f0f: y = 16'h200;
			16'h5f10: y = 16'h200;
			16'h5f11: y = 16'h200;
			16'h5f12: y = 16'h200;
			16'h5f13: y = 16'h200;
			16'h5f14: y = 16'h200;
			16'h5f15: y = 16'h200;
			16'h5f16: y = 16'h200;
			16'h5f17: y = 16'h200;
			16'h5f18: y = 16'h200;
			16'h5f19: y = 16'h200;
			16'h5f1a: y = 16'h200;
			16'h5f1b: y = 16'h200;
			16'h5f1c: y = 16'h200;
			16'h5f1d: y = 16'h200;
			16'h5f1e: y = 16'h200;
			16'h5f1f: y = 16'h200;
			16'h5f20: y = 16'h200;
			16'h5f21: y = 16'h200;
			16'h5f22: y = 16'h200;
			16'h5f23: y = 16'h200;
			16'h5f24: y = 16'h200;
			16'h5f25: y = 16'h200;
			16'h5f26: y = 16'h200;
			16'h5f27: y = 16'h200;
			16'h5f28: y = 16'h200;
			16'h5f29: y = 16'h200;
			16'h5f2a: y = 16'h200;
			16'h5f2b: y = 16'h200;
			16'h5f2c: y = 16'h200;
			16'h5f2d: y = 16'h200;
			16'h5f2e: y = 16'h200;
			16'h5f2f: y = 16'h200;
			16'h5f30: y = 16'h200;
			16'h5f31: y = 16'h200;
			16'h5f32: y = 16'h200;
			16'h5f33: y = 16'h200;
			16'h5f34: y = 16'h200;
			16'h5f35: y = 16'h200;
			16'h5f36: y = 16'h200;
			16'h5f37: y = 16'h200;
			16'h5f38: y = 16'h200;
			16'h5f39: y = 16'h200;
			16'h5f3a: y = 16'h200;
			16'h5f3b: y = 16'h200;
			16'h5f3c: y = 16'h200;
			16'h5f3d: y = 16'h200;
			16'h5f3e: y = 16'h200;
			16'h5f3f: y = 16'h200;
			16'h5f40: y = 16'h200;
			16'h5f41: y = 16'h200;
			16'h5f42: y = 16'h200;
			16'h5f43: y = 16'h200;
			16'h5f44: y = 16'h200;
			16'h5f45: y = 16'h200;
			16'h5f46: y = 16'h200;
			16'h5f47: y = 16'h200;
			16'h5f48: y = 16'h200;
			16'h5f49: y = 16'h200;
			16'h5f4a: y = 16'h200;
			16'h5f4b: y = 16'h200;
			16'h5f4c: y = 16'h200;
			16'h5f4d: y = 16'h200;
			16'h5f4e: y = 16'h200;
			16'h5f4f: y = 16'h200;
			16'h5f50: y = 16'h200;
			16'h5f51: y = 16'h200;
			16'h5f52: y = 16'h200;
			16'h5f53: y = 16'h200;
			16'h5f54: y = 16'h200;
			16'h5f55: y = 16'h200;
			16'h5f56: y = 16'h200;
			16'h5f57: y = 16'h200;
			16'h5f58: y = 16'h200;
			16'h5f59: y = 16'h200;
			16'h5f5a: y = 16'h200;
			16'h5f5b: y = 16'h200;
			16'h5f5c: y = 16'h200;
			16'h5f5d: y = 16'h200;
			16'h5f5e: y = 16'h200;
			16'h5f5f: y = 16'h200;
			16'h5f60: y = 16'h200;
			16'h5f61: y = 16'h200;
			16'h5f62: y = 16'h200;
			16'h5f63: y = 16'h200;
			16'h5f64: y = 16'h200;
			16'h5f65: y = 16'h200;
			16'h5f66: y = 16'h200;
			16'h5f67: y = 16'h200;
			16'h5f68: y = 16'h200;
			16'h5f69: y = 16'h200;
			16'h5f6a: y = 16'h200;
			16'h5f6b: y = 16'h200;
			16'h5f6c: y = 16'h200;
			16'h5f6d: y = 16'h200;
			16'h5f6e: y = 16'h200;
			16'h5f6f: y = 16'h200;
			16'h5f70: y = 16'h200;
			16'h5f71: y = 16'h200;
			16'h5f72: y = 16'h200;
			16'h5f73: y = 16'h200;
			16'h5f74: y = 16'h200;
			16'h5f75: y = 16'h200;
			16'h5f76: y = 16'h200;
			16'h5f77: y = 16'h200;
			16'h5f78: y = 16'h200;
			16'h5f79: y = 16'h200;
			16'h5f7a: y = 16'h200;
			16'h5f7b: y = 16'h200;
			16'h5f7c: y = 16'h200;
			16'h5f7d: y = 16'h200;
			16'h5f7e: y = 16'h200;
			16'h5f7f: y = 16'h200;
			16'h5f80: y = 16'h200;
			16'h5f81: y = 16'h200;
			16'h5f82: y = 16'h200;
			16'h5f83: y = 16'h200;
			16'h5f84: y = 16'h200;
			16'h5f85: y = 16'h200;
			16'h5f86: y = 16'h200;
			16'h5f87: y = 16'h200;
			16'h5f88: y = 16'h200;
			16'h5f89: y = 16'h200;
			16'h5f8a: y = 16'h200;
			16'h5f8b: y = 16'h200;
			16'h5f8c: y = 16'h200;
			16'h5f8d: y = 16'h200;
			16'h5f8e: y = 16'h200;
			16'h5f8f: y = 16'h200;
			16'h5f90: y = 16'h200;
			16'h5f91: y = 16'h200;
			16'h5f92: y = 16'h200;
			16'h5f93: y = 16'h200;
			16'h5f94: y = 16'h200;
			16'h5f95: y = 16'h200;
			16'h5f96: y = 16'h200;
			16'h5f97: y = 16'h200;
			16'h5f98: y = 16'h200;
			16'h5f99: y = 16'h200;
			16'h5f9a: y = 16'h200;
			16'h5f9b: y = 16'h200;
			16'h5f9c: y = 16'h200;
			16'h5f9d: y = 16'h200;
			16'h5f9e: y = 16'h200;
			16'h5f9f: y = 16'h200;
			16'h5fa0: y = 16'h200;
			16'h5fa1: y = 16'h200;
			16'h5fa2: y = 16'h200;
			16'h5fa3: y = 16'h200;
			16'h5fa4: y = 16'h200;
			16'h5fa5: y = 16'h200;
			16'h5fa6: y = 16'h200;
			16'h5fa7: y = 16'h200;
			16'h5fa8: y = 16'h200;
			16'h5fa9: y = 16'h200;
			16'h5faa: y = 16'h200;
			16'h5fab: y = 16'h200;
			16'h5fac: y = 16'h200;
			16'h5fad: y = 16'h200;
			16'h5fae: y = 16'h200;
			16'h5faf: y = 16'h200;
			16'h5fb0: y = 16'h200;
			16'h5fb1: y = 16'h200;
			16'h5fb2: y = 16'h200;
			16'h5fb3: y = 16'h200;
			16'h5fb4: y = 16'h200;
			16'h5fb5: y = 16'h200;
			16'h5fb6: y = 16'h200;
			16'h5fb7: y = 16'h200;
			16'h5fb8: y = 16'h200;
			16'h5fb9: y = 16'h200;
			16'h5fba: y = 16'h200;
			16'h5fbb: y = 16'h200;
			16'h5fbc: y = 16'h200;
			16'h5fbd: y = 16'h200;
			16'h5fbe: y = 16'h200;
			16'h5fbf: y = 16'h200;
			16'h5fc0: y = 16'h200;
			16'h5fc1: y = 16'h200;
			16'h5fc2: y = 16'h200;
			16'h5fc3: y = 16'h200;
			16'h5fc4: y = 16'h200;
			16'h5fc5: y = 16'h200;
			16'h5fc6: y = 16'h200;
			16'h5fc7: y = 16'h200;
			16'h5fc8: y = 16'h200;
			16'h5fc9: y = 16'h200;
			16'h5fca: y = 16'h200;
			16'h5fcb: y = 16'h200;
			16'h5fcc: y = 16'h200;
			16'h5fcd: y = 16'h200;
			16'h5fce: y = 16'h200;
			16'h5fcf: y = 16'h200;
			16'h5fd0: y = 16'h200;
			16'h5fd1: y = 16'h200;
			16'h5fd2: y = 16'h200;
			16'h5fd3: y = 16'h200;
			16'h5fd4: y = 16'h200;
			16'h5fd5: y = 16'h200;
			16'h5fd6: y = 16'h200;
			16'h5fd7: y = 16'h200;
			16'h5fd8: y = 16'h200;
			16'h5fd9: y = 16'h200;
			16'h5fda: y = 16'h200;
			16'h5fdb: y = 16'h200;
			16'h5fdc: y = 16'h200;
			16'h5fdd: y = 16'h200;
			16'h5fde: y = 16'h200;
			16'h5fdf: y = 16'h200;
			16'h5fe0: y = 16'h200;
			16'h5fe1: y = 16'h200;
			16'h5fe2: y = 16'h200;
			16'h5fe3: y = 16'h200;
			16'h5fe4: y = 16'h200;
			16'h5fe5: y = 16'h200;
			16'h5fe6: y = 16'h200;
			16'h5fe7: y = 16'h200;
			16'h5fe8: y = 16'h200;
			16'h5fe9: y = 16'h200;
			16'h5fea: y = 16'h200;
			16'h5feb: y = 16'h200;
			16'h5fec: y = 16'h200;
			16'h5fed: y = 16'h200;
			16'h5fee: y = 16'h200;
			16'h5fef: y = 16'h200;
			16'h5ff0: y = 16'h200;
			16'h5ff1: y = 16'h200;
			16'h5ff2: y = 16'h200;
			16'h5ff3: y = 16'h200;
			16'h5ff4: y = 16'h200;
			16'h5ff5: y = 16'h200;
			16'h5ff6: y = 16'h200;
			16'h5ff7: y = 16'h200;
			16'h5ff8: y = 16'h200;
			16'h5ff9: y = 16'h200;
			16'h5ffa: y = 16'h200;
			16'h5ffb: y = 16'h200;
			16'h5ffc: y = 16'h200;
			16'h5ffd: y = 16'h200;
			16'h5ffe: y = 16'h200;
			16'h5fff: y = 16'h200;
			16'h6000: y = 16'h200;
			16'h6001: y = 16'h200;
			16'h6002: y = 16'h200;
			16'h6003: y = 16'h200;
			16'h6004: y = 16'h200;
			16'h6005: y = 16'h200;
			16'h6006: y = 16'h200;
			16'h6007: y = 16'h200;
			16'h6008: y = 16'h200;
			16'h6009: y = 16'h200;
			16'h600a: y = 16'h200;
			16'h600b: y = 16'h200;
			16'h600c: y = 16'h200;
			16'h600d: y = 16'h200;
			16'h600e: y = 16'h200;
			16'h600f: y = 16'h200;
			16'h6010: y = 16'h200;
			16'h6011: y = 16'h200;
			16'h6012: y = 16'h200;
			16'h6013: y = 16'h200;
			16'h6014: y = 16'h200;
			16'h6015: y = 16'h200;
			16'h6016: y = 16'h200;
			16'h6017: y = 16'h200;
			16'h6018: y = 16'h200;
			16'h6019: y = 16'h200;
			16'h601a: y = 16'h200;
			16'h601b: y = 16'h200;
			16'h601c: y = 16'h200;
			16'h601d: y = 16'h200;
			16'h601e: y = 16'h200;
			16'h601f: y = 16'h200;
			16'h6020: y = 16'h200;
			16'h6021: y = 16'h200;
			16'h6022: y = 16'h200;
			16'h6023: y = 16'h200;
			16'h6024: y = 16'h200;
			16'h6025: y = 16'h200;
			16'h6026: y = 16'h200;
			16'h6027: y = 16'h200;
			16'h6028: y = 16'h200;
			16'h6029: y = 16'h200;
			16'h602a: y = 16'h200;
			16'h602b: y = 16'h200;
			16'h602c: y = 16'h200;
			16'h602d: y = 16'h200;
			16'h602e: y = 16'h200;
			16'h602f: y = 16'h200;
			16'h6030: y = 16'h200;
			16'h6031: y = 16'h200;
			16'h6032: y = 16'h200;
			16'h6033: y = 16'h200;
			16'h6034: y = 16'h200;
			16'h6035: y = 16'h200;
			16'h6036: y = 16'h200;
			16'h6037: y = 16'h200;
			16'h6038: y = 16'h200;
			16'h6039: y = 16'h200;
			16'h603a: y = 16'h200;
			16'h603b: y = 16'h200;
			16'h603c: y = 16'h200;
			16'h603d: y = 16'h200;
			16'h603e: y = 16'h200;
			16'h603f: y = 16'h200;
			16'h6040: y = 16'h200;
			16'h6041: y = 16'h200;
			16'h6042: y = 16'h200;
			16'h6043: y = 16'h200;
			16'h6044: y = 16'h200;
			16'h6045: y = 16'h200;
			16'h6046: y = 16'h200;
			16'h6047: y = 16'h200;
			16'h6048: y = 16'h200;
			16'h6049: y = 16'h200;
			16'h604a: y = 16'h200;
			16'h604b: y = 16'h200;
			16'h604c: y = 16'h200;
			16'h604d: y = 16'h200;
			16'h604e: y = 16'h200;
			16'h604f: y = 16'h200;
			16'h6050: y = 16'h200;
			16'h6051: y = 16'h200;
			16'h6052: y = 16'h200;
			16'h6053: y = 16'h200;
			16'h6054: y = 16'h200;
			16'h6055: y = 16'h200;
			16'h6056: y = 16'h200;
			16'h6057: y = 16'h200;
			16'h6058: y = 16'h200;
			16'h6059: y = 16'h200;
			16'h605a: y = 16'h200;
			16'h605b: y = 16'h200;
			16'h605c: y = 16'h200;
			16'h605d: y = 16'h200;
			16'h605e: y = 16'h200;
			16'h605f: y = 16'h200;
			16'h6060: y = 16'h200;
			16'h6061: y = 16'h200;
			16'h6062: y = 16'h200;
			16'h6063: y = 16'h200;
			16'h6064: y = 16'h200;
			16'h6065: y = 16'h200;
			16'h6066: y = 16'h200;
			16'h6067: y = 16'h200;
			16'h6068: y = 16'h200;
			16'h6069: y = 16'h200;
			16'h606a: y = 16'h200;
			16'h606b: y = 16'h200;
			16'h606c: y = 16'h200;
			16'h606d: y = 16'h200;
			16'h606e: y = 16'h200;
			16'h606f: y = 16'h200;
			16'h6070: y = 16'h200;
			16'h6071: y = 16'h200;
			16'h6072: y = 16'h200;
			16'h6073: y = 16'h200;
			16'h6074: y = 16'h200;
			16'h6075: y = 16'h200;
			16'h6076: y = 16'h200;
			16'h6077: y = 16'h200;
			16'h6078: y = 16'h200;
			16'h6079: y = 16'h200;
			16'h607a: y = 16'h200;
			16'h607b: y = 16'h200;
			16'h607c: y = 16'h200;
			16'h607d: y = 16'h200;
			16'h607e: y = 16'h200;
			16'h607f: y = 16'h200;
			16'h6080: y = 16'h200;
			16'h6081: y = 16'h200;
			16'h6082: y = 16'h200;
			16'h6083: y = 16'h200;
			16'h6084: y = 16'h200;
			16'h6085: y = 16'h200;
			16'h6086: y = 16'h200;
			16'h6087: y = 16'h200;
			16'h6088: y = 16'h200;
			16'h6089: y = 16'h200;
			16'h608a: y = 16'h200;
			16'h608b: y = 16'h200;
			16'h608c: y = 16'h200;
			16'h608d: y = 16'h200;
			16'h608e: y = 16'h200;
			16'h608f: y = 16'h200;
			16'h6090: y = 16'h200;
			16'h6091: y = 16'h200;
			16'h6092: y = 16'h200;
			16'h6093: y = 16'h200;
			16'h6094: y = 16'h200;
			16'h6095: y = 16'h200;
			16'h6096: y = 16'h200;
			16'h6097: y = 16'h200;
			16'h6098: y = 16'h200;
			16'h6099: y = 16'h200;
			16'h609a: y = 16'h200;
			16'h609b: y = 16'h200;
			16'h609c: y = 16'h200;
			16'h609d: y = 16'h200;
			16'h609e: y = 16'h200;
			16'h609f: y = 16'h200;
			16'h60a0: y = 16'h200;
			16'h60a1: y = 16'h200;
			16'h60a2: y = 16'h200;
			16'h60a3: y = 16'h200;
			16'h60a4: y = 16'h200;
			16'h60a5: y = 16'h200;
			16'h60a6: y = 16'h200;
			16'h60a7: y = 16'h200;
			16'h60a8: y = 16'h200;
			16'h60a9: y = 16'h200;
			16'h60aa: y = 16'h200;
			16'h60ab: y = 16'h200;
			16'h60ac: y = 16'h200;
			16'h60ad: y = 16'h200;
			16'h60ae: y = 16'h200;
			16'h60af: y = 16'h200;
			16'h60b0: y = 16'h200;
			16'h60b1: y = 16'h200;
			16'h60b2: y = 16'h200;
			16'h60b3: y = 16'h200;
			16'h60b4: y = 16'h200;
			16'h60b5: y = 16'h200;
			16'h60b6: y = 16'h200;
			16'h60b7: y = 16'h200;
			16'h60b8: y = 16'h200;
			16'h60b9: y = 16'h200;
			16'h60ba: y = 16'h200;
			16'h60bb: y = 16'h200;
			16'h60bc: y = 16'h200;
			16'h60bd: y = 16'h200;
			16'h60be: y = 16'h200;
			16'h60bf: y = 16'h200;
			16'h60c0: y = 16'h200;
			16'h60c1: y = 16'h200;
			16'h60c2: y = 16'h200;
			16'h60c3: y = 16'h200;
			16'h60c4: y = 16'h200;
			16'h60c5: y = 16'h200;
			16'h60c6: y = 16'h200;
			16'h60c7: y = 16'h200;
			16'h60c8: y = 16'h200;
			16'h60c9: y = 16'h200;
			16'h60ca: y = 16'h200;
			16'h60cb: y = 16'h200;
			16'h60cc: y = 16'h200;
			16'h60cd: y = 16'h200;
			16'h60ce: y = 16'h200;
			16'h60cf: y = 16'h200;
			16'h60d0: y = 16'h200;
			16'h60d1: y = 16'h200;
			16'h60d2: y = 16'h200;
			16'h60d3: y = 16'h200;
			16'h60d4: y = 16'h200;
			16'h60d5: y = 16'h200;
			16'h60d6: y = 16'h200;
			16'h60d7: y = 16'h200;
			16'h60d8: y = 16'h200;
			16'h60d9: y = 16'h200;
			16'h60da: y = 16'h200;
			16'h60db: y = 16'h200;
			16'h60dc: y = 16'h200;
			16'h60dd: y = 16'h200;
			16'h60de: y = 16'h200;
			16'h60df: y = 16'h200;
			16'h60e0: y = 16'h200;
			16'h60e1: y = 16'h200;
			16'h60e2: y = 16'h200;
			16'h60e3: y = 16'h200;
			16'h60e4: y = 16'h200;
			16'h60e5: y = 16'h200;
			16'h60e6: y = 16'h200;
			16'h60e7: y = 16'h200;
			16'h60e8: y = 16'h200;
			16'h60e9: y = 16'h200;
			16'h60ea: y = 16'h200;
			16'h60eb: y = 16'h200;
			16'h60ec: y = 16'h200;
			16'h60ed: y = 16'h200;
			16'h60ee: y = 16'h200;
			16'h60ef: y = 16'h200;
			16'h60f0: y = 16'h200;
			16'h60f1: y = 16'h200;
			16'h60f2: y = 16'h200;
			16'h60f3: y = 16'h200;
			16'h60f4: y = 16'h200;
			16'h60f5: y = 16'h200;
			16'h60f6: y = 16'h200;
			16'h60f7: y = 16'h200;
			16'h60f8: y = 16'h200;
			16'h60f9: y = 16'h200;
			16'h60fa: y = 16'h200;
			16'h60fb: y = 16'h200;
			16'h60fc: y = 16'h200;
			16'h60fd: y = 16'h200;
			16'h60fe: y = 16'h200;
			16'h60ff: y = 16'h200;
			16'h6100: y = 16'h200;
			16'h6101: y = 16'h200;
			16'h6102: y = 16'h200;
			16'h6103: y = 16'h200;
			16'h6104: y = 16'h200;
			16'h6105: y = 16'h200;
			16'h6106: y = 16'h200;
			16'h6107: y = 16'h200;
			16'h6108: y = 16'h200;
			16'h6109: y = 16'h200;
			16'h610a: y = 16'h200;
			16'h610b: y = 16'h200;
			16'h610c: y = 16'h200;
			16'h610d: y = 16'h200;
			16'h610e: y = 16'h200;
			16'h610f: y = 16'h200;
			16'h6110: y = 16'h200;
			16'h6111: y = 16'h200;
			16'h6112: y = 16'h200;
			16'h6113: y = 16'h200;
			16'h6114: y = 16'h200;
			16'h6115: y = 16'h200;
			16'h6116: y = 16'h200;
			16'h6117: y = 16'h200;
			16'h6118: y = 16'h200;
			16'h6119: y = 16'h200;
			16'h611a: y = 16'h200;
			16'h611b: y = 16'h200;
			16'h611c: y = 16'h200;
			16'h611d: y = 16'h200;
			16'h611e: y = 16'h200;
			16'h611f: y = 16'h200;
			16'h6120: y = 16'h200;
			16'h6121: y = 16'h200;
			16'h6122: y = 16'h200;
			16'h6123: y = 16'h200;
			16'h6124: y = 16'h200;
			16'h6125: y = 16'h200;
			16'h6126: y = 16'h200;
			16'h6127: y = 16'h200;
			16'h6128: y = 16'h200;
			16'h6129: y = 16'h200;
			16'h612a: y = 16'h200;
			16'h612b: y = 16'h200;
			16'h612c: y = 16'h200;
			16'h612d: y = 16'h200;
			16'h612e: y = 16'h200;
			16'h612f: y = 16'h200;
			16'h6130: y = 16'h200;
			16'h6131: y = 16'h200;
			16'h6132: y = 16'h200;
			16'h6133: y = 16'h200;
			16'h6134: y = 16'h200;
			16'h6135: y = 16'h200;
			16'h6136: y = 16'h200;
			16'h6137: y = 16'h200;
			16'h6138: y = 16'h200;
			16'h6139: y = 16'h200;
			16'h613a: y = 16'h200;
			16'h613b: y = 16'h200;
			16'h613c: y = 16'h200;
			16'h613d: y = 16'h200;
			16'h613e: y = 16'h200;
			16'h613f: y = 16'h200;
			16'h6140: y = 16'h200;
			16'h6141: y = 16'h200;
			16'h6142: y = 16'h200;
			16'h6143: y = 16'h200;
			16'h6144: y = 16'h200;
			16'h6145: y = 16'h200;
			16'h6146: y = 16'h200;
			16'h6147: y = 16'h200;
			16'h6148: y = 16'h200;
			16'h6149: y = 16'h200;
			16'h614a: y = 16'h200;
			16'h614b: y = 16'h200;
			16'h614c: y = 16'h200;
			16'h614d: y = 16'h200;
			16'h614e: y = 16'h200;
			16'h614f: y = 16'h200;
			16'h6150: y = 16'h200;
			16'h6151: y = 16'h200;
			16'h6152: y = 16'h200;
			16'h6153: y = 16'h200;
			16'h6154: y = 16'h200;
			16'h6155: y = 16'h200;
			16'h6156: y = 16'h200;
			16'h6157: y = 16'h200;
			16'h6158: y = 16'h200;
			16'h6159: y = 16'h200;
			16'h615a: y = 16'h200;
			16'h615b: y = 16'h200;
			16'h615c: y = 16'h200;
			16'h615d: y = 16'h200;
			16'h615e: y = 16'h200;
			16'h615f: y = 16'h200;
			16'h6160: y = 16'h200;
			16'h6161: y = 16'h200;
			16'h6162: y = 16'h200;
			16'h6163: y = 16'h200;
			16'h6164: y = 16'h200;
			16'h6165: y = 16'h200;
			16'h6166: y = 16'h200;
			16'h6167: y = 16'h200;
			16'h6168: y = 16'h200;
			16'h6169: y = 16'h200;
			16'h616a: y = 16'h200;
			16'h616b: y = 16'h200;
			16'h616c: y = 16'h200;
			16'h616d: y = 16'h200;
			16'h616e: y = 16'h200;
			16'h616f: y = 16'h200;
			16'h6170: y = 16'h200;
			16'h6171: y = 16'h200;
			16'h6172: y = 16'h200;
			16'h6173: y = 16'h200;
			16'h6174: y = 16'h200;
			16'h6175: y = 16'h200;
			16'h6176: y = 16'h200;
			16'h6177: y = 16'h200;
			16'h6178: y = 16'h200;
			16'h6179: y = 16'h200;
			16'h617a: y = 16'h200;
			16'h617b: y = 16'h200;
			16'h617c: y = 16'h200;
			16'h617d: y = 16'h200;
			16'h617e: y = 16'h200;
			16'h617f: y = 16'h200;
			16'h6180: y = 16'h200;
			16'h6181: y = 16'h200;
			16'h6182: y = 16'h200;
			16'h6183: y = 16'h200;
			16'h6184: y = 16'h200;
			16'h6185: y = 16'h200;
			16'h6186: y = 16'h200;
			16'h6187: y = 16'h200;
			16'h6188: y = 16'h200;
			16'h6189: y = 16'h200;
			16'h618a: y = 16'h200;
			16'h618b: y = 16'h200;
			16'h618c: y = 16'h200;
			16'h618d: y = 16'h200;
			16'h618e: y = 16'h200;
			16'h618f: y = 16'h200;
			16'h6190: y = 16'h200;
			16'h6191: y = 16'h200;
			16'h6192: y = 16'h200;
			16'h6193: y = 16'h200;
			16'h6194: y = 16'h200;
			16'h6195: y = 16'h200;
			16'h6196: y = 16'h200;
			16'h6197: y = 16'h200;
			16'h6198: y = 16'h200;
			16'h6199: y = 16'h200;
			16'h619a: y = 16'h200;
			16'h619b: y = 16'h200;
			16'h619c: y = 16'h200;
			16'h619d: y = 16'h200;
			16'h619e: y = 16'h200;
			16'h619f: y = 16'h200;
			16'h61a0: y = 16'h200;
			16'h61a1: y = 16'h200;
			16'h61a2: y = 16'h200;
			16'h61a3: y = 16'h200;
			16'h61a4: y = 16'h200;
			16'h61a5: y = 16'h200;
			16'h61a6: y = 16'h200;
			16'h61a7: y = 16'h200;
			16'h61a8: y = 16'h200;
			16'h61a9: y = 16'h200;
			16'h61aa: y = 16'h200;
			16'h61ab: y = 16'h200;
			16'h61ac: y = 16'h200;
			16'h61ad: y = 16'h200;
			16'h61ae: y = 16'h200;
			16'h61af: y = 16'h200;
			16'h61b0: y = 16'h200;
			16'h61b1: y = 16'h200;
			16'h61b2: y = 16'h200;
			16'h61b3: y = 16'h200;
			16'h61b4: y = 16'h200;
			16'h61b5: y = 16'h200;
			16'h61b6: y = 16'h200;
			16'h61b7: y = 16'h200;
			16'h61b8: y = 16'h200;
			16'h61b9: y = 16'h200;
			16'h61ba: y = 16'h200;
			16'h61bb: y = 16'h200;
			16'h61bc: y = 16'h200;
			16'h61bd: y = 16'h200;
			16'h61be: y = 16'h200;
			16'h61bf: y = 16'h200;
			16'h61c0: y = 16'h200;
			16'h61c1: y = 16'h200;
			16'h61c2: y = 16'h200;
			16'h61c3: y = 16'h200;
			16'h61c4: y = 16'h200;
			16'h61c5: y = 16'h200;
			16'h61c6: y = 16'h200;
			16'h61c7: y = 16'h200;
			16'h61c8: y = 16'h200;
			16'h61c9: y = 16'h200;
			16'h61ca: y = 16'h200;
			16'h61cb: y = 16'h200;
			16'h61cc: y = 16'h200;
			16'h61cd: y = 16'h200;
			16'h61ce: y = 16'h200;
			16'h61cf: y = 16'h200;
			16'h61d0: y = 16'h200;
			16'h61d1: y = 16'h200;
			16'h61d2: y = 16'h200;
			16'h61d3: y = 16'h200;
			16'h61d4: y = 16'h200;
			16'h61d5: y = 16'h200;
			16'h61d6: y = 16'h200;
			16'h61d7: y = 16'h200;
			16'h61d8: y = 16'h200;
			16'h61d9: y = 16'h200;
			16'h61da: y = 16'h200;
			16'h61db: y = 16'h200;
			16'h61dc: y = 16'h200;
			16'h61dd: y = 16'h200;
			16'h61de: y = 16'h200;
			16'h61df: y = 16'h200;
			16'h61e0: y = 16'h200;
			16'h61e1: y = 16'h200;
			16'h61e2: y = 16'h200;
			16'h61e3: y = 16'h200;
			16'h61e4: y = 16'h200;
			16'h61e5: y = 16'h200;
			16'h61e6: y = 16'h200;
			16'h61e7: y = 16'h200;
			16'h61e8: y = 16'h200;
			16'h61e9: y = 16'h200;
			16'h61ea: y = 16'h200;
			16'h61eb: y = 16'h200;
			16'h61ec: y = 16'h200;
			16'h61ed: y = 16'h200;
			16'h61ee: y = 16'h200;
			16'h61ef: y = 16'h200;
			16'h61f0: y = 16'h200;
			16'h61f1: y = 16'h200;
			16'h61f2: y = 16'h200;
			16'h61f3: y = 16'h200;
			16'h61f4: y = 16'h200;
			16'h61f5: y = 16'h200;
			16'h61f6: y = 16'h200;
			16'h61f7: y = 16'h200;
			16'h61f8: y = 16'h200;
			16'h61f9: y = 16'h200;
			16'h61fa: y = 16'h200;
			16'h61fb: y = 16'h200;
			16'h61fc: y = 16'h200;
			16'h61fd: y = 16'h200;
			16'h61fe: y = 16'h200;
			16'h61ff: y = 16'h200;
			16'h6200: y = 16'h200;
			16'h6201: y = 16'h200;
			16'h6202: y = 16'h200;
			16'h6203: y = 16'h200;
			16'h6204: y = 16'h200;
			16'h6205: y = 16'h200;
			16'h6206: y = 16'h200;
			16'h6207: y = 16'h200;
			16'h6208: y = 16'h200;
			16'h6209: y = 16'h200;
			16'h620a: y = 16'h200;
			16'h620b: y = 16'h200;
			16'h620c: y = 16'h200;
			16'h620d: y = 16'h200;
			16'h620e: y = 16'h200;
			16'h620f: y = 16'h200;
			16'h6210: y = 16'h200;
			16'h6211: y = 16'h200;
			16'h6212: y = 16'h200;
			16'h6213: y = 16'h200;
			16'h6214: y = 16'h200;
			16'h6215: y = 16'h200;
			16'h6216: y = 16'h200;
			16'h6217: y = 16'h200;
			16'h6218: y = 16'h200;
			16'h6219: y = 16'h200;
			16'h621a: y = 16'h200;
			16'h621b: y = 16'h200;
			16'h621c: y = 16'h200;
			16'h621d: y = 16'h200;
			16'h621e: y = 16'h200;
			16'h621f: y = 16'h200;
			16'h6220: y = 16'h200;
			16'h6221: y = 16'h200;
			16'h6222: y = 16'h200;
			16'h6223: y = 16'h200;
			16'h6224: y = 16'h200;
			16'h6225: y = 16'h200;
			16'h6226: y = 16'h200;
			16'h6227: y = 16'h200;
			16'h6228: y = 16'h200;
			16'h6229: y = 16'h200;
			16'h622a: y = 16'h200;
			16'h622b: y = 16'h200;
			16'h622c: y = 16'h200;
			16'h622d: y = 16'h200;
			16'h622e: y = 16'h200;
			16'h622f: y = 16'h200;
			16'h6230: y = 16'h200;
			16'h6231: y = 16'h200;
			16'h6232: y = 16'h200;
			16'h6233: y = 16'h200;
			16'h6234: y = 16'h200;
			16'h6235: y = 16'h200;
			16'h6236: y = 16'h200;
			16'h6237: y = 16'h200;
			16'h6238: y = 16'h200;
			16'h6239: y = 16'h200;
			16'h623a: y = 16'h200;
			16'h623b: y = 16'h200;
			16'h623c: y = 16'h200;
			16'h623d: y = 16'h200;
			16'h623e: y = 16'h200;
			16'h623f: y = 16'h200;
			16'h6240: y = 16'h200;
			16'h6241: y = 16'h200;
			16'h6242: y = 16'h200;
			16'h6243: y = 16'h200;
			16'h6244: y = 16'h200;
			16'h6245: y = 16'h200;
			16'h6246: y = 16'h200;
			16'h6247: y = 16'h200;
			16'h6248: y = 16'h200;
			16'h6249: y = 16'h200;
			16'h624a: y = 16'h200;
			16'h624b: y = 16'h200;
			16'h624c: y = 16'h200;
			16'h624d: y = 16'h200;
			16'h624e: y = 16'h200;
			16'h624f: y = 16'h200;
			16'h6250: y = 16'h200;
			16'h6251: y = 16'h200;
			16'h6252: y = 16'h200;
			16'h6253: y = 16'h200;
			16'h6254: y = 16'h200;
			16'h6255: y = 16'h200;
			16'h6256: y = 16'h200;
			16'h6257: y = 16'h200;
			16'h6258: y = 16'h200;
			16'h6259: y = 16'h200;
			16'h625a: y = 16'h200;
			16'h625b: y = 16'h200;
			16'h625c: y = 16'h200;
			16'h625d: y = 16'h200;
			16'h625e: y = 16'h200;
			16'h625f: y = 16'h200;
			16'h6260: y = 16'h200;
			16'h6261: y = 16'h200;
			16'h6262: y = 16'h200;
			16'h6263: y = 16'h200;
			16'h6264: y = 16'h200;
			16'h6265: y = 16'h200;
			16'h6266: y = 16'h200;
			16'h6267: y = 16'h200;
			16'h6268: y = 16'h200;
			16'h6269: y = 16'h200;
			16'h626a: y = 16'h200;
			16'h626b: y = 16'h200;
			16'h626c: y = 16'h200;
			16'h626d: y = 16'h200;
			16'h626e: y = 16'h200;
			16'h626f: y = 16'h200;
			16'h6270: y = 16'h200;
			16'h6271: y = 16'h200;
			16'h6272: y = 16'h200;
			16'h6273: y = 16'h200;
			16'h6274: y = 16'h200;
			16'h6275: y = 16'h200;
			16'h6276: y = 16'h200;
			16'h6277: y = 16'h200;
			16'h6278: y = 16'h200;
			16'h6279: y = 16'h200;
			16'h627a: y = 16'h200;
			16'h627b: y = 16'h200;
			16'h627c: y = 16'h200;
			16'h627d: y = 16'h200;
			16'h627e: y = 16'h200;
			16'h627f: y = 16'h200;
			16'h6280: y = 16'h200;
			16'h6281: y = 16'h200;
			16'h6282: y = 16'h200;
			16'h6283: y = 16'h200;
			16'h6284: y = 16'h200;
			16'h6285: y = 16'h200;
			16'h6286: y = 16'h200;
			16'h6287: y = 16'h200;
			16'h6288: y = 16'h200;
			16'h6289: y = 16'h200;
			16'h628a: y = 16'h200;
			16'h628b: y = 16'h200;
			16'h628c: y = 16'h200;
			16'h628d: y = 16'h200;
			16'h628e: y = 16'h200;
			16'h628f: y = 16'h200;
			16'h6290: y = 16'h200;
			16'h6291: y = 16'h200;
			16'h6292: y = 16'h200;
			16'h6293: y = 16'h200;
			16'h6294: y = 16'h200;
			16'h6295: y = 16'h200;
			16'h6296: y = 16'h200;
			16'h6297: y = 16'h200;
			16'h6298: y = 16'h200;
			16'h6299: y = 16'h200;
			16'h629a: y = 16'h200;
			16'h629b: y = 16'h200;
			16'h629c: y = 16'h200;
			16'h629d: y = 16'h200;
			16'h629e: y = 16'h200;
			16'h629f: y = 16'h200;
			16'h62a0: y = 16'h200;
			16'h62a1: y = 16'h200;
			16'h62a2: y = 16'h200;
			16'h62a3: y = 16'h200;
			16'h62a4: y = 16'h200;
			16'h62a5: y = 16'h200;
			16'h62a6: y = 16'h200;
			16'h62a7: y = 16'h200;
			16'h62a8: y = 16'h200;
			16'h62a9: y = 16'h200;
			16'h62aa: y = 16'h200;
			16'h62ab: y = 16'h200;
			16'h62ac: y = 16'h200;
			16'h62ad: y = 16'h200;
			16'h62ae: y = 16'h200;
			16'h62af: y = 16'h200;
			16'h62b0: y = 16'h200;
			16'h62b1: y = 16'h200;
			16'h62b2: y = 16'h200;
			16'h62b3: y = 16'h200;
			16'h62b4: y = 16'h200;
			16'h62b5: y = 16'h200;
			16'h62b6: y = 16'h200;
			16'h62b7: y = 16'h200;
			16'h62b8: y = 16'h200;
			16'h62b9: y = 16'h200;
			16'h62ba: y = 16'h200;
			16'h62bb: y = 16'h200;
			16'h62bc: y = 16'h200;
			16'h62bd: y = 16'h200;
			16'h62be: y = 16'h200;
			16'h62bf: y = 16'h200;
			16'h62c0: y = 16'h200;
			16'h62c1: y = 16'h200;
			16'h62c2: y = 16'h200;
			16'h62c3: y = 16'h200;
			16'h62c4: y = 16'h200;
			16'h62c5: y = 16'h200;
			16'h62c6: y = 16'h200;
			16'h62c7: y = 16'h200;
			16'h62c8: y = 16'h200;
			16'h62c9: y = 16'h200;
			16'h62ca: y = 16'h200;
			16'h62cb: y = 16'h200;
			16'h62cc: y = 16'h200;
			16'h62cd: y = 16'h200;
			16'h62ce: y = 16'h200;
			16'h62cf: y = 16'h200;
			16'h62d0: y = 16'h200;
			16'h62d1: y = 16'h200;
			16'h62d2: y = 16'h200;
			16'h62d3: y = 16'h200;
			16'h62d4: y = 16'h200;
			16'h62d5: y = 16'h200;
			16'h62d6: y = 16'h200;
			16'h62d7: y = 16'h200;
			16'h62d8: y = 16'h200;
			16'h62d9: y = 16'h200;
			16'h62da: y = 16'h200;
			16'h62db: y = 16'h200;
			16'h62dc: y = 16'h200;
			16'h62dd: y = 16'h200;
			16'h62de: y = 16'h200;
			16'h62df: y = 16'h200;
			16'h62e0: y = 16'h200;
			16'h62e1: y = 16'h200;
			16'h62e2: y = 16'h200;
			16'h62e3: y = 16'h200;
			16'h62e4: y = 16'h200;
			16'h62e5: y = 16'h200;
			16'h62e6: y = 16'h200;
			16'h62e7: y = 16'h200;
			16'h62e8: y = 16'h200;
			16'h62e9: y = 16'h200;
			16'h62ea: y = 16'h200;
			16'h62eb: y = 16'h200;
			16'h62ec: y = 16'h200;
			16'h62ed: y = 16'h200;
			16'h62ee: y = 16'h200;
			16'h62ef: y = 16'h200;
			16'h62f0: y = 16'h200;
			16'h62f1: y = 16'h200;
			16'h62f2: y = 16'h200;
			16'h62f3: y = 16'h200;
			16'h62f4: y = 16'h200;
			16'h62f5: y = 16'h200;
			16'h62f6: y = 16'h200;
			16'h62f7: y = 16'h200;
			16'h62f8: y = 16'h200;
			16'h62f9: y = 16'h200;
			16'h62fa: y = 16'h200;
			16'h62fb: y = 16'h200;
			16'h62fc: y = 16'h200;
			16'h62fd: y = 16'h200;
			16'h62fe: y = 16'h200;
			16'h62ff: y = 16'h200;
			16'h6300: y = 16'h200;
			16'h6301: y = 16'h200;
			16'h6302: y = 16'h200;
			16'h6303: y = 16'h200;
			16'h6304: y = 16'h200;
			16'h6305: y = 16'h200;
			16'h6306: y = 16'h200;
			16'h6307: y = 16'h200;
			16'h6308: y = 16'h200;
			16'h6309: y = 16'h200;
			16'h630a: y = 16'h200;
			16'h630b: y = 16'h200;
			16'h630c: y = 16'h200;
			16'h630d: y = 16'h200;
			16'h630e: y = 16'h200;
			16'h630f: y = 16'h200;
			16'h6310: y = 16'h200;
			16'h6311: y = 16'h200;
			16'h6312: y = 16'h200;
			16'h6313: y = 16'h200;
			16'h6314: y = 16'h200;
			16'h6315: y = 16'h200;
			16'h6316: y = 16'h200;
			16'h6317: y = 16'h200;
			16'h6318: y = 16'h200;
			16'h6319: y = 16'h200;
			16'h631a: y = 16'h200;
			16'h631b: y = 16'h200;
			16'h631c: y = 16'h200;
			16'h631d: y = 16'h200;
			16'h631e: y = 16'h200;
			16'h631f: y = 16'h200;
			16'h6320: y = 16'h200;
			16'h6321: y = 16'h200;
			16'h6322: y = 16'h200;
			16'h6323: y = 16'h200;
			16'h6324: y = 16'h200;
			16'h6325: y = 16'h200;
			16'h6326: y = 16'h200;
			16'h6327: y = 16'h200;
			16'h6328: y = 16'h200;
			16'h6329: y = 16'h200;
			16'h632a: y = 16'h200;
			16'h632b: y = 16'h200;
			16'h632c: y = 16'h200;
			16'h632d: y = 16'h200;
			16'h632e: y = 16'h200;
			16'h632f: y = 16'h200;
			16'h6330: y = 16'h200;
			16'h6331: y = 16'h200;
			16'h6332: y = 16'h200;
			16'h6333: y = 16'h200;
			16'h6334: y = 16'h200;
			16'h6335: y = 16'h200;
			16'h6336: y = 16'h200;
			16'h6337: y = 16'h200;
			16'h6338: y = 16'h200;
			16'h6339: y = 16'h200;
			16'h633a: y = 16'h200;
			16'h633b: y = 16'h200;
			16'h633c: y = 16'h200;
			16'h633d: y = 16'h200;
			16'h633e: y = 16'h200;
			16'h633f: y = 16'h200;
			16'h6340: y = 16'h200;
			16'h6341: y = 16'h200;
			16'h6342: y = 16'h200;
			16'h6343: y = 16'h200;
			16'h6344: y = 16'h200;
			16'h6345: y = 16'h200;
			16'h6346: y = 16'h200;
			16'h6347: y = 16'h200;
			16'h6348: y = 16'h200;
			16'h6349: y = 16'h200;
			16'h634a: y = 16'h200;
			16'h634b: y = 16'h200;
			16'h634c: y = 16'h200;
			16'h634d: y = 16'h200;
			16'h634e: y = 16'h200;
			16'h634f: y = 16'h200;
			16'h6350: y = 16'h200;
			16'h6351: y = 16'h200;
			16'h6352: y = 16'h200;
			16'h6353: y = 16'h200;
			16'h6354: y = 16'h200;
			16'h6355: y = 16'h200;
			16'h6356: y = 16'h200;
			16'h6357: y = 16'h200;
			16'h6358: y = 16'h200;
			16'h6359: y = 16'h200;
			16'h635a: y = 16'h200;
			16'h635b: y = 16'h200;
			16'h635c: y = 16'h200;
			16'h635d: y = 16'h200;
			16'h635e: y = 16'h200;
			16'h635f: y = 16'h200;
			16'h6360: y = 16'h200;
			16'h6361: y = 16'h200;
			16'h6362: y = 16'h200;
			16'h6363: y = 16'h200;
			16'h6364: y = 16'h200;
			16'h6365: y = 16'h200;
			16'h6366: y = 16'h200;
			16'h6367: y = 16'h200;
			16'h6368: y = 16'h200;
			16'h6369: y = 16'h200;
			16'h636a: y = 16'h200;
			16'h636b: y = 16'h200;
			16'h636c: y = 16'h200;
			16'h636d: y = 16'h200;
			16'h636e: y = 16'h200;
			16'h636f: y = 16'h200;
			16'h6370: y = 16'h200;
			16'h6371: y = 16'h200;
			16'h6372: y = 16'h200;
			16'h6373: y = 16'h200;
			16'h6374: y = 16'h200;
			16'h6375: y = 16'h200;
			16'h6376: y = 16'h200;
			16'h6377: y = 16'h200;
			16'h6378: y = 16'h200;
			16'h6379: y = 16'h200;
			16'h637a: y = 16'h200;
			16'h637b: y = 16'h200;
			16'h637c: y = 16'h200;
			16'h637d: y = 16'h200;
			16'h637e: y = 16'h200;
			16'h637f: y = 16'h200;
			16'h6380: y = 16'h200;
			16'h6381: y = 16'h200;
			16'h6382: y = 16'h200;
			16'h6383: y = 16'h200;
			16'h6384: y = 16'h200;
			16'h6385: y = 16'h200;
			16'h6386: y = 16'h200;
			16'h6387: y = 16'h200;
			16'h6388: y = 16'h200;
			16'h6389: y = 16'h200;
			16'h638a: y = 16'h200;
			16'h638b: y = 16'h200;
			16'h638c: y = 16'h200;
			16'h638d: y = 16'h200;
			16'h638e: y = 16'h200;
			16'h638f: y = 16'h200;
			16'h6390: y = 16'h200;
			16'h6391: y = 16'h200;
			16'h6392: y = 16'h200;
			16'h6393: y = 16'h200;
			16'h6394: y = 16'h200;
			16'h6395: y = 16'h200;
			16'h6396: y = 16'h200;
			16'h6397: y = 16'h200;
			16'h6398: y = 16'h200;
			16'h6399: y = 16'h200;
			16'h639a: y = 16'h200;
			16'h639b: y = 16'h200;
			16'h639c: y = 16'h200;
			16'h639d: y = 16'h200;
			16'h639e: y = 16'h200;
			16'h639f: y = 16'h200;
			16'h63a0: y = 16'h200;
			16'h63a1: y = 16'h200;
			16'h63a2: y = 16'h200;
			16'h63a3: y = 16'h200;
			16'h63a4: y = 16'h200;
			16'h63a5: y = 16'h200;
			16'h63a6: y = 16'h200;
			16'h63a7: y = 16'h200;
			16'h63a8: y = 16'h200;
			16'h63a9: y = 16'h200;
			16'h63aa: y = 16'h200;
			16'h63ab: y = 16'h200;
			16'h63ac: y = 16'h200;
			16'h63ad: y = 16'h200;
			16'h63ae: y = 16'h200;
			16'h63af: y = 16'h200;
			16'h63b0: y = 16'h200;
			16'h63b1: y = 16'h200;
			16'h63b2: y = 16'h200;
			16'h63b3: y = 16'h200;
			16'h63b4: y = 16'h200;
			16'h63b5: y = 16'h200;
			16'h63b6: y = 16'h200;
			16'h63b7: y = 16'h200;
			16'h63b8: y = 16'h200;
			16'h63b9: y = 16'h200;
			16'h63ba: y = 16'h200;
			16'h63bb: y = 16'h200;
			16'h63bc: y = 16'h200;
			16'h63bd: y = 16'h200;
			16'h63be: y = 16'h200;
			16'h63bf: y = 16'h200;
			16'h63c0: y = 16'h200;
			16'h63c1: y = 16'h200;
			16'h63c2: y = 16'h200;
			16'h63c3: y = 16'h200;
			16'h63c4: y = 16'h200;
			16'h63c5: y = 16'h200;
			16'h63c6: y = 16'h200;
			16'h63c7: y = 16'h200;
			16'h63c8: y = 16'h200;
			16'h63c9: y = 16'h200;
			16'h63ca: y = 16'h200;
			16'h63cb: y = 16'h200;
			16'h63cc: y = 16'h200;
			16'h63cd: y = 16'h200;
			16'h63ce: y = 16'h200;
			16'h63cf: y = 16'h200;
			16'h63d0: y = 16'h200;
			16'h63d1: y = 16'h200;
			16'h63d2: y = 16'h200;
			16'h63d3: y = 16'h200;
			16'h63d4: y = 16'h200;
			16'h63d5: y = 16'h200;
			16'h63d6: y = 16'h200;
			16'h63d7: y = 16'h200;
			16'h63d8: y = 16'h200;
			16'h63d9: y = 16'h200;
			16'h63da: y = 16'h200;
			16'h63db: y = 16'h200;
			16'h63dc: y = 16'h200;
			16'h63dd: y = 16'h200;
			16'h63de: y = 16'h200;
			16'h63df: y = 16'h200;
			16'h63e0: y = 16'h200;
			16'h63e1: y = 16'h200;
			16'h63e2: y = 16'h200;
			16'h63e3: y = 16'h200;
			16'h63e4: y = 16'h200;
			16'h63e5: y = 16'h200;
			16'h63e6: y = 16'h200;
			16'h63e7: y = 16'h200;
			16'h63e8: y = 16'h200;
			16'h63e9: y = 16'h200;
			16'h63ea: y = 16'h200;
			16'h63eb: y = 16'h200;
			16'h63ec: y = 16'h200;
			16'h63ed: y = 16'h200;
			16'h63ee: y = 16'h200;
			16'h63ef: y = 16'h200;
			16'h63f0: y = 16'h200;
			16'h63f1: y = 16'h200;
			16'h63f2: y = 16'h200;
			16'h63f3: y = 16'h200;
			16'h63f4: y = 16'h200;
			16'h63f5: y = 16'h200;
			16'h63f6: y = 16'h200;
			16'h63f7: y = 16'h200;
			16'h63f8: y = 16'h200;
			16'h63f9: y = 16'h200;
			16'h63fa: y = 16'h200;
			16'h63fb: y = 16'h200;
			16'h63fc: y = 16'h200;
			16'h63fd: y = 16'h200;
			16'h63fe: y = 16'h200;
			16'h63ff: y = 16'h200;
			16'h6400: y = 16'h200;
			16'h6401: y = 16'h200;
			16'h6402: y = 16'h200;
			16'h6403: y = 16'h200;
			16'h6404: y = 16'h200;
			16'h6405: y = 16'h200;
			16'h6406: y = 16'h200;
			16'h6407: y = 16'h200;
			16'h6408: y = 16'h200;
			16'h6409: y = 16'h200;
			16'h640a: y = 16'h200;
			16'h640b: y = 16'h200;
			16'h640c: y = 16'h200;
			16'h640d: y = 16'h200;
			16'h640e: y = 16'h200;
			16'h640f: y = 16'h200;
			16'h6410: y = 16'h200;
			16'h6411: y = 16'h200;
			16'h6412: y = 16'h200;
			16'h6413: y = 16'h200;
			16'h6414: y = 16'h200;
			16'h6415: y = 16'h200;
			16'h6416: y = 16'h200;
			16'h6417: y = 16'h200;
			16'h6418: y = 16'h200;
			16'h6419: y = 16'h200;
			16'h641a: y = 16'h200;
			16'h641b: y = 16'h200;
			16'h641c: y = 16'h200;
			16'h641d: y = 16'h200;
			16'h641e: y = 16'h200;
			16'h641f: y = 16'h200;
			16'h6420: y = 16'h200;
			16'h6421: y = 16'h200;
			16'h6422: y = 16'h200;
			16'h6423: y = 16'h200;
			16'h6424: y = 16'h200;
			16'h6425: y = 16'h200;
			16'h6426: y = 16'h200;
			16'h6427: y = 16'h200;
			16'h6428: y = 16'h200;
			16'h6429: y = 16'h200;
			16'h642a: y = 16'h200;
			16'h642b: y = 16'h200;
			16'h642c: y = 16'h200;
			16'h642d: y = 16'h200;
			16'h642e: y = 16'h200;
			16'h642f: y = 16'h200;
			16'h6430: y = 16'h200;
			16'h6431: y = 16'h200;
			16'h6432: y = 16'h200;
			16'h6433: y = 16'h200;
			16'h6434: y = 16'h200;
			16'h6435: y = 16'h200;
			16'h6436: y = 16'h200;
			16'h6437: y = 16'h200;
			16'h6438: y = 16'h200;
			16'h6439: y = 16'h200;
			16'h643a: y = 16'h200;
			16'h643b: y = 16'h200;
			16'h643c: y = 16'h200;
			16'h643d: y = 16'h200;
			16'h643e: y = 16'h200;
			16'h643f: y = 16'h200;
			16'h6440: y = 16'h200;
			16'h6441: y = 16'h200;
			16'h6442: y = 16'h200;
			16'h6443: y = 16'h200;
			16'h6444: y = 16'h200;
			16'h6445: y = 16'h200;
			16'h6446: y = 16'h200;
			16'h6447: y = 16'h200;
			16'h6448: y = 16'h200;
			16'h6449: y = 16'h200;
			16'h644a: y = 16'h200;
			16'h644b: y = 16'h200;
			16'h644c: y = 16'h200;
			16'h644d: y = 16'h200;
			16'h644e: y = 16'h200;
			16'h644f: y = 16'h200;
			16'h6450: y = 16'h200;
			16'h6451: y = 16'h200;
			16'h6452: y = 16'h200;
			16'h6453: y = 16'h200;
			16'h6454: y = 16'h200;
			16'h6455: y = 16'h200;
			16'h6456: y = 16'h200;
			16'h6457: y = 16'h200;
			16'h6458: y = 16'h200;
			16'h6459: y = 16'h200;
			16'h645a: y = 16'h200;
			16'h645b: y = 16'h200;
			16'h645c: y = 16'h200;
			16'h645d: y = 16'h200;
			16'h645e: y = 16'h200;
			16'h645f: y = 16'h200;
			16'h6460: y = 16'h200;
			16'h6461: y = 16'h200;
			16'h6462: y = 16'h200;
			16'h6463: y = 16'h200;
			16'h6464: y = 16'h200;
			16'h6465: y = 16'h200;
			16'h6466: y = 16'h200;
			16'h6467: y = 16'h200;
			16'h6468: y = 16'h200;
			16'h6469: y = 16'h200;
			16'h646a: y = 16'h200;
			16'h646b: y = 16'h200;
			16'h646c: y = 16'h200;
			16'h646d: y = 16'h200;
			16'h646e: y = 16'h200;
			16'h646f: y = 16'h200;
			16'h6470: y = 16'h200;
			16'h6471: y = 16'h200;
			16'h6472: y = 16'h200;
			16'h6473: y = 16'h200;
			16'h6474: y = 16'h200;
			16'h6475: y = 16'h200;
			16'h6476: y = 16'h200;
			16'h6477: y = 16'h200;
			16'h6478: y = 16'h200;
			16'h6479: y = 16'h200;
			16'h647a: y = 16'h200;
			16'h647b: y = 16'h200;
			16'h647c: y = 16'h200;
			16'h647d: y = 16'h200;
			16'h647e: y = 16'h200;
			16'h647f: y = 16'h200;
			16'h6480: y = 16'h200;
			16'h6481: y = 16'h200;
			16'h6482: y = 16'h200;
			16'h6483: y = 16'h200;
			16'h6484: y = 16'h200;
			16'h6485: y = 16'h200;
			16'h6486: y = 16'h200;
			16'h6487: y = 16'h200;
			16'h6488: y = 16'h200;
			16'h6489: y = 16'h200;
			16'h648a: y = 16'h200;
			16'h648b: y = 16'h200;
			16'h648c: y = 16'h200;
			16'h648d: y = 16'h200;
			16'h648e: y = 16'h200;
			16'h648f: y = 16'h200;
			16'h6490: y = 16'h200;
			16'h6491: y = 16'h200;
			16'h6492: y = 16'h200;
			16'h6493: y = 16'h200;
			16'h6494: y = 16'h200;
			16'h6495: y = 16'h200;
			16'h6496: y = 16'h200;
			16'h6497: y = 16'h200;
			16'h6498: y = 16'h200;
			16'h6499: y = 16'h200;
			16'h649a: y = 16'h200;
			16'h649b: y = 16'h200;
			16'h649c: y = 16'h200;
			16'h649d: y = 16'h200;
			16'h649e: y = 16'h200;
			16'h649f: y = 16'h200;
			16'h64a0: y = 16'h200;
			16'h64a1: y = 16'h200;
			16'h64a2: y = 16'h200;
			16'h64a3: y = 16'h200;
			16'h64a4: y = 16'h200;
			16'h64a5: y = 16'h200;
			16'h64a6: y = 16'h200;
			16'h64a7: y = 16'h200;
			16'h64a8: y = 16'h200;
			16'h64a9: y = 16'h200;
			16'h64aa: y = 16'h200;
			16'h64ab: y = 16'h200;
			16'h64ac: y = 16'h200;
			16'h64ad: y = 16'h200;
			16'h64ae: y = 16'h200;
			16'h64af: y = 16'h200;
			16'h64b0: y = 16'h200;
			16'h64b1: y = 16'h200;
			16'h64b2: y = 16'h200;
			16'h64b3: y = 16'h200;
			16'h64b4: y = 16'h200;
			16'h64b5: y = 16'h200;
			16'h64b6: y = 16'h200;
			16'h64b7: y = 16'h200;
			16'h64b8: y = 16'h200;
			16'h64b9: y = 16'h200;
			16'h64ba: y = 16'h200;
			16'h64bb: y = 16'h200;
			16'h64bc: y = 16'h200;
			16'h64bd: y = 16'h200;
			16'h64be: y = 16'h200;
			16'h64bf: y = 16'h200;
			16'h64c0: y = 16'h200;
			16'h64c1: y = 16'h200;
			16'h64c2: y = 16'h200;
			16'h64c3: y = 16'h200;
			16'h64c4: y = 16'h200;
			16'h64c5: y = 16'h200;
			16'h64c6: y = 16'h200;
			16'h64c7: y = 16'h200;
			16'h64c8: y = 16'h200;
			16'h64c9: y = 16'h200;
			16'h64ca: y = 16'h200;
			16'h64cb: y = 16'h200;
			16'h64cc: y = 16'h200;
			16'h64cd: y = 16'h200;
			16'h64ce: y = 16'h200;
			16'h64cf: y = 16'h200;
			16'h64d0: y = 16'h200;
			16'h64d1: y = 16'h200;
			16'h64d2: y = 16'h200;
			16'h64d3: y = 16'h200;
			16'h64d4: y = 16'h200;
			16'h64d5: y = 16'h200;
			16'h64d6: y = 16'h200;
			16'h64d7: y = 16'h200;
			16'h64d8: y = 16'h200;
			16'h64d9: y = 16'h200;
			16'h64da: y = 16'h200;
			16'h64db: y = 16'h200;
			16'h64dc: y = 16'h200;
			16'h64dd: y = 16'h200;
			16'h64de: y = 16'h200;
			16'h64df: y = 16'h200;
			16'h64e0: y = 16'h200;
			16'h64e1: y = 16'h200;
			16'h64e2: y = 16'h200;
			16'h64e3: y = 16'h200;
			16'h64e4: y = 16'h200;
			16'h64e5: y = 16'h200;
			16'h64e6: y = 16'h200;
			16'h64e7: y = 16'h200;
			16'h64e8: y = 16'h200;
			16'h64e9: y = 16'h200;
			16'h64ea: y = 16'h200;
			16'h64eb: y = 16'h200;
			16'h64ec: y = 16'h200;
			16'h64ed: y = 16'h200;
			16'h64ee: y = 16'h200;
			16'h64ef: y = 16'h200;
			16'h64f0: y = 16'h200;
			16'h64f1: y = 16'h200;
			16'h64f2: y = 16'h200;
			16'h64f3: y = 16'h200;
			16'h64f4: y = 16'h200;
			16'h64f5: y = 16'h200;
			16'h64f6: y = 16'h200;
			16'h64f7: y = 16'h200;
			16'h64f8: y = 16'h200;
			16'h64f9: y = 16'h200;
			16'h64fa: y = 16'h200;
			16'h64fb: y = 16'h200;
			16'h64fc: y = 16'h200;
			16'h64fd: y = 16'h200;
			16'h64fe: y = 16'h200;
			16'h64ff: y = 16'h200;
			16'h6500: y = 16'h200;
			16'h6501: y = 16'h200;
			16'h6502: y = 16'h200;
			16'h6503: y = 16'h200;
			16'h6504: y = 16'h200;
			16'h6505: y = 16'h200;
			16'h6506: y = 16'h200;
			16'h6507: y = 16'h200;
			16'h6508: y = 16'h200;
			16'h6509: y = 16'h200;
			16'h650a: y = 16'h200;
			16'h650b: y = 16'h200;
			16'h650c: y = 16'h200;
			16'h650d: y = 16'h200;
			16'h650e: y = 16'h200;
			16'h650f: y = 16'h200;
			16'h6510: y = 16'h200;
			16'h6511: y = 16'h200;
			16'h6512: y = 16'h200;
			16'h6513: y = 16'h200;
			16'h6514: y = 16'h200;
			16'h6515: y = 16'h200;
			16'h6516: y = 16'h200;
			16'h6517: y = 16'h200;
			16'h6518: y = 16'h200;
			16'h6519: y = 16'h200;
			16'h651a: y = 16'h200;
			16'h651b: y = 16'h200;
			16'h651c: y = 16'h200;
			16'h651d: y = 16'h200;
			16'h651e: y = 16'h200;
			16'h651f: y = 16'h200;
			16'h6520: y = 16'h200;
			16'h6521: y = 16'h200;
			16'h6522: y = 16'h200;
			16'h6523: y = 16'h200;
			16'h6524: y = 16'h200;
			16'h6525: y = 16'h200;
			16'h6526: y = 16'h200;
			16'h6527: y = 16'h200;
			16'h6528: y = 16'h200;
			16'h6529: y = 16'h200;
			16'h652a: y = 16'h200;
			16'h652b: y = 16'h200;
			16'h652c: y = 16'h200;
			16'h652d: y = 16'h200;
			16'h652e: y = 16'h200;
			16'h652f: y = 16'h200;
			16'h6530: y = 16'h200;
			16'h6531: y = 16'h200;
			16'h6532: y = 16'h200;
			16'h6533: y = 16'h200;
			16'h6534: y = 16'h200;
			16'h6535: y = 16'h200;
			16'h6536: y = 16'h200;
			16'h6537: y = 16'h200;
			16'h6538: y = 16'h200;
			16'h6539: y = 16'h200;
			16'h653a: y = 16'h200;
			16'h653b: y = 16'h200;
			16'h653c: y = 16'h200;
			16'h653d: y = 16'h200;
			16'h653e: y = 16'h200;
			16'h653f: y = 16'h200;
			16'h6540: y = 16'h200;
			16'h6541: y = 16'h200;
			16'h6542: y = 16'h200;
			16'h6543: y = 16'h200;
			16'h6544: y = 16'h200;
			16'h6545: y = 16'h200;
			16'h6546: y = 16'h200;
			16'h6547: y = 16'h200;
			16'h6548: y = 16'h200;
			16'h6549: y = 16'h200;
			16'h654a: y = 16'h200;
			16'h654b: y = 16'h200;
			16'h654c: y = 16'h200;
			16'h654d: y = 16'h200;
			16'h654e: y = 16'h200;
			16'h654f: y = 16'h200;
			16'h6550: y = 16'h200;
			16'h6551: y = 16'h200;
			16'h6552: y = 16'h200;
			16'h6553: y = 16'h200;
			16'h6554: y = 16'h200;
			16'h6555: y = 16'h200;
			16'h6556: y = 16'h200;
			16'h6557: y = 16'h200;
			16'h6558: y = 16'h200;
			16'h6559: y = 16'h200;
			16'h655a: y = 16'h200;
			16'h655b: y = 16'h200;
			16'h655c: y = 16'h200;
			16'h655d: y = 16'h200;
			16'h655e: y = 16'h200;
			16'h655f: y = 16'h200;
			16'h6560: y = 16'h200;
			16'h6561: y = 16'h200;
			16'h6562: y = 16'h200;
			16'h6563: y = 16'h200;
			16'h6564: y = 16'h200;
			16'h6565: y = 16'h200;
			16'h6566: y = 16'h200;
			16'h6567: y = 16'h200;
			16'h6568: y = 16'h200;
			16'h6569: y = 16'h200;
			16'h656a: y = 16'h200;
			16'h656b: y = 16'h200;
			16'h656c: y = 16'h200;
			16'h656d: y = 16'h200;
			16'h656e: y = 16'h200;
			16'h656f: y = 16'h200;
			16'h6570: y = 16'h200;
			16'h6571: y = 16'h200;
			16'h6572: y = 16'h200;
			16'h6573: y = 16'h200;
			16'h6574: y = 16'h200;
			16'h6575: y = 16'h200;
			16'h6576: y = 16'h200;
			16'h6577: y = 16'h200;
			16'h6578: y = 16'h200;
			16'h6579: y = 16'h200;
			16'h657a: y = 16'h200;
			16'h657b: y = 16'h200;
			16'h657c: y = 16'h200;
			16'h657d: y = 16'h200;
			16'h657e: y = 16'h200;
			16'h657f: y = 16'h200;
			16'h6580: y = 16'h200;
			16'h6581: y = 16'h200;
			16'h6582: y = 16'h200;
			16'h6583: y = 16'h200;
			16'h6584: y = 16'h200;
			16'h6585: y = 16'h200;
			16'h6586: y = 16'h200;
			16'h6587: y = 16'h200;
			16'h6588: y = 16'h200;
			16'h6589: y = 16'h200;
			16'h658a: y = 16'h200;
			16'h658b: y = 16'h200;
			16'h658c: y = 16'h200;
			16'h658d: y = 16'h200;
			16'h658e: y = 16'h200;
			16'h658f: y = 16'h200;
			16'h6590: y = 16'h200;
			16'h6591: y = 16'h200;
			16'h6592: y = 16'h200;
			16'h6593: y = 16'h200;
			16'h6594: y = 16'h200;
			16'h6595: y = 16'h200;
			16'h6596: y = 16'h200;
			16'h6597: y = 16'h200;
			16'h6598: y = 16'h200;
			16'h6599: y = 16'h200;
			16'h659a: y = 16'h200;
			16'h659b: y = 16'h200;
			16'h659c: y = 16'h200;
			16'h659d: y = 16'h200;
			16'h659e: y = 16'h200;
			16'h659f: y = 16'h200;
			16'h65a0: y = 16'h200;
			16'h65a1: y = 16'h200;
			16'h65a2: y = 16'h200;
			16'h65a3: y = 16'h200;
			16'h65a4: y = 16'h200;
			16'h65a5: y = 16'h200;
			16'h65a6: y = 16'h200;
			16'h65a7: y = 16'h200;
			16'h65a8: y = 16'h200;
			16'h65a9: y = 16'h200;
			16'h65aa: y = 16'h200;
			16'h65ab: y = 16'h200;
			16'h65ac: y = 16'h200;
			16'h65ad: y = 16'h200;
			16'h65ae: y = 16'h200;
			16'h65af: y = 16'h200;
			16'h65b0: y = 16'h200;
			16'h65b1: y = 16'h200;
			16'h65b2: y = 16'h200;
			16'h65b3: y = 16'h200;
			16'h65b4: y = 16'h200;
			16'h65b5: y = 16'h200;
			16'h65b6: y = 16'h200;
			16'h65b7: y = 16'h200;
			16'h65b8: y = 16'h200;
			16'h65b9: y = 16'h200;
			16'h65ba: y = 16'h200;
			16'h65bb: y = 16'h200;
			16'h65bc: y = 16'h200;
			16'h65bd: y = 16'h200;
			16'h65be: y = 16'h200;
			16'h65bf: y = 16'h200;
			16'h65c0: y = 16'h200;
			16'h65c1: y = 16'h200;
			16'h65c2: y = 16'h200;
			16'h65c3: y = 16'h200;
			16'h65c4: y = 16'h200;
			16'h65c5: y = 16'h200;
			16'h65c6: y = 16'h200;
			16'h65c7: y = 16'h200;
			16'h65c8: y = 16'h200;
			16'h65c9: y = 16'h200;
			16'h65ca: y = 16'h200;
			16'h65cb: y = 16'h200;
			16'h65cc: y = 16'h200;
			16'h65cd: y = 16'h200;
			16'h65ce: y = 16'h200;
			16'h65cf: y = 16'h200;
			16'h65d0: y = 16'h200;
			16'h65d1: y = 16'h200;
			16'h65d2: y = 16'h200;
			16'h65d3: y = 16'h200;
			16'h65d4: y = 16'h200;
			16'h65d5: y = 16'h200;
			16'h65d6: y = 16'h200;
			16'h65d7: y = 16'h200;
			16'h65d8: y = 16'h200;
			16'h65d9: y = 16'h200;
			16'h65da: y = 16'h200;
			16'h65db: y = 16'h200;
			16'h65dc: y = 16'h200;
			16'h65dd: y = 16'h200;
			16'h65de: y = 16'h200;
			16'h65df: y = 16'h200;
			16'h65e0: y = 16'h200;
			16'h65e1: y = 16'h200;
			16'h65e2: y = 16'h200;
			16'h65e3: y = 16'h200;
			16'h65e4: y = 16'h200;
			16'h65e5: y = 16'h200;
			16'h65e6: y = 16'h200;
			16'h65e7: y = 16'h200;
			16'h65e8: y = 16'h200;
			16'h65e9: y = 16'h200;
			16'h65ea: y = 16'h200;
			16'h65eb: y = 16'h200;
			16'h65ec: y = 16'h200;
			16'h65ed: y = 16'h200;
			16'h65ee: y = 16'h200;
			16'h65ef: y = 16'h200;
			16'h65f0: y = 16'h200;
			16'h65f1: y = 16'h200;
			16'h65f2: y = 16'h200;
			16'h65f3: y = 16'h200;
			16'h65f4: y = 16'h200;
			16'h65f5: y = 16'h200;
			16'h65f6: y = 16'h200;
			16'h65f7: y = 16'h200;
			16'h65f8: y = 16'h200;
			16'h65f9: y = 16'h200;
			16'h65fa: y = 16'h200;
			16'h65fb: y = 16'h200;
			16'h65fc: y = 16'h200;
			16'h65fd: y = 16'h200;
			16'h65fe: y = 16'h200;
			16'h65ff: y = 16'h200;
			16'h6600: y = 16'h200;
			16'h6601: y = 16'h200;
			16'h6602: y = 16'h200;
			16'h6603: y = 16'h200;
			16'h6604: y = 16'h200;
			16'h6605: y = 16'h200;
			16'h6606: y = 16'h200;
			16'h6607: y = 16'h200;
			16'h6608: y = 16'h200;
			16'h6609: y = 16'h200;
			16'h660a: y = 16'h200;
			16'h660b: y = 16'h200;
			16'h660c: y = 16'h200;
			16'h660d: y = 16'h200;
			16'h660e: y = 16'h200;
			16'h660f: y = 16'h200;
			16'h6610: y = 16'h200;
			16'h6611: y = 16'h200;
			16'h6612: y = 16'h200;
			16'h6613: y = 16'h200;
			16'h6614: y = 16'h200;
			16'h6615: y = 16'h200;
			16'h6616: y = 16'h200;
			16'h6617: y = 16'h200;
			16'h6618: y = 16'h200;
			16'h6619: y = 16'h200;
			16'h661a: y = 16'h200;
			16'h661b: y = 16'h200;
			16'h661c: y = 16'h200;
			16'h661d: y = 16'h200;
			16'h661e: y = 16'h200;
			16'h661f: y = 16'h200;
			16'h6620: y = 16'h200;
			16'h6621: y = 16'h200;
			16'h6622: y = 16'h200;
			16'h6623: y = 16'h200;
			16'h6624: y = 16'h200;
			16'h6625: y = 16'h200;
			16'h6626: y = 16'h200;
			16'h6627: y = 16'h200;
			16'h6628: y = 16'h200;
			16'h6629: y = 16'h200;
			16'h662a: y = 16'h200;
			16'h662b: y = 16'h200;
			16'h662c: y = 16'h200;
			16'h662d: y = 16'h200;
			16'h662e: y = 16'h200;
			16'h662f: y = 16'h200;
			16'h6630: y = 16'h200;
			16'h6631: y = 16'h200;
			16'h6632: y = 16'h200;
			16'h6633: y = 16'h200;
			16'h6634: y = 16'h200;
			16'h6635: y = 16'h200;
			16'h6636: y = 16'h200;
			16'h6637: y = 16'h200;
			16'h6638: y = 16'h200;
			16'h6639: y = 16'h200;
			16'h663a: y = 16'h200;
			16'h663b: y = 16'h200;
			16'h663c: y = 16'h200;
			16'h663d: y = 16'h200;
			16'h663e: y = 16'h200;
			16'h663f: y = 16'h200;
			16'h6640: y = 16'h200;
			16'h6641: y = 16'h200;
			16'h6642: y = 16'h200;
			16'h6643: y = 16'h200;
			16'h6644: y = 16'h200;
			16'h6645: y = 16'h200;
			16'h6646: y = 16'h200;
			16'h6647: y = 16'h200;
			16'h6648: y = 16'h200;
			16'h6649: y = 16'h200;
			16'h664a: y = 16'h200;
			16'h664b: y = 16'h200;
			16'h664c: y = 16'h200;
			16'h664d: y = 16'h200;
			16'h664e: y = 16'h200;
			16'h664f: y = 16'h200;
			16'h6650: y = 16'h200;
			16'h6651: y = 16'h200;
			16'h6652: y = 16'h200;
			16'h6653: y = 16'h200;
			16'h6654: y = 16'h200;
			16'h6655: y = 16'h200;
			16'h6656: y = 16'h200;
			16'h6657: y = 16'h200;
			16'h6658: y = 16'h200;
			16'h6659: y = 16'h200;
			16'h665a: y = 16'h200;
			16'h665b: y = 16'h200;
			16'h665c: y = 16'h200;
			16'h665d: y = 16'h200;
			16'h665e: y = 16'h200;
			16'h665f: y = 16'h200;
			16'h6660: y = 16'h200;
			16'h6661: y = 16'h200;
			16'h6662: y = 16'h200;
			16'h6663: y = 16'h200;
			16'h6664: y = 16'h200;
			16'h6665: y = 16'h200;
			16'h6666: y = 16'h200;
			16'h6667: y = 16'h200;
			16'h6668: y = 16'h200;
			16'h6669: y = 16'h200;
			16'h666a: y = 16'h200;
			16'h666b: y = 16'h200;
			16'h666c: y = 16'h200;
			16'h666d: y = 16'h200;
			16'h666e: y = 16'h200;
			16'h666f: y = 16'h200;
			16'h6670: y = 16'h200;
			16'h6671: y = 16'h200;
			16'h6672: y = 16'h200;
			16'h6673: y = 16'h200;
			16'h6674: y = 16'h200;
			16'h6675: y = 16'h200;
			16'h6676: y = 16'h200;
			16'h6677: y = 16'h200;
			16'h6678: y = 16'h200;
			16'h6679: y = 16'h200;
			16'h667a: y = 16'h200;
			16'h667b: y = 16'h200;
			16'h667c: y = 16'h200;
			16'h667d: y = 16'h200;
			16'h667e: y = 16'h200;
			16'h667f: y = 16'h200;
			16'h6680: y = 16'h200;
			16'h6681: y = 16'h200;
			16'h6682: y = 16'h200;
			16'h6683: y = 16'h200;
			16'h6684: y = 16'h200;
			16'h6685: y = 16'h200;
			16'h6686: y = 16'h200;
			16'h6687: y = 16'h200;
			16'h6688: y = 16'h200;
			16'h6689: y = 16'h200;
			16'h668a: y = 16'h200;
			16'h668b: y = 16'h200;
			16'h668c: y = 16'h200;
			16'h668d: y = 16'h200;
			16'h668e: y = 16'h200;
			16'h668f: y = 16'h200;
			16'h6690: y = 16'h200;
			16'h6691: y = 16'h200;
			16'h6692: y = 16'h200;
			16'h6693: y = 16'h200;
			16'h6694: y = 16'h200;
			16'h6695: y = 16'h200;
			16'h6696: y = 16'h200;
			16'h6697: y = 16'h200;
			16'h6698: y = 16'h200;
			16'h6699: y = 16'h200;
			16'h669a: y = 16'h200;
			16'h669b: y = 16'h200;
			16'h669c: y = 16'h200;
			16'h669d: y = 16'h200;
			16'h669e: y = 16'h200;
			16'h669f: y = 16'h200;
			16'h66a0: y = 16'h200;
			16'h66a1: y = 16'h200;
			16'h66a2: y = 16'h200;
			16'h66a3: y = 16'h200;
			16'h66a4: y = 16'h200;
			16'h66a5: y = 16'h200;
			16'h66a6: y = 16'h200;
			16'h66a7: y = 16'h200;
			16'h66a8: y = 16'h200;
			16'h66a9: y = 16'h200;
			16'h66aa: y = 16'h200;
			16'h66ab: y = 16'h200;
			16'h66ac: y = 16'h200;
			16'h66ad: y = 16'h200;
			16'h66ae: y = 16'h200;
			16'h66af: y = 16'h200;
			16'h66b0: y = 16'h200;
			16'h66b1: y = 16'h200;
			16'h66b2: y = 16'h200;
			16'h66b3: y = 16'h200;
			16'h66b4: y = 16'h200;
			16'h66b5: y = 16'h200;
			16'h66b6: y = 16'h200;
			16'h66b7: y = 16'h200;
			16'h66b8: y = 16'h200;
			16'h66b9: y = 16'h200;
			16'h66ba: y = 16'h200;
			16'h66bb: y = 16'h200;
			16'h66bc: y = 16'h200;
			16'h66bd: y = 16'h200;
			16'h66be: y = 16'h200;
			16'h66bf: y = 16'h200;
			16'h66c0: y = 16'h200;
			16'h66c1: y = 16'h200;
			16'h66c2: y = 16'h200;
			16'h66c3: y = 16'h200;
			16'h66c4: y = 16'h200;
			16'h66c5: y = 16'h200;
			16'h66c6: y = 16'h200;
			16'h66c7: y = 16'h200;
			16'h66c8: y = 16'h200;
			16'h66c9: y = 16'h200;
			16'h66ca: y = 16'h200;
			16'h66cb: y = 16'h200;
			16'h66cc: y = 16'h200;
			16'h66cd: y = 16'h200;
			16'h66ce: y = 16'h200;
			16'h66cf: y = 16'h200;
			16'h66d0: y = 16'h200;
			16'h66d1: y = 16'h200;
			16'h66d2: y = 16'h200;
			16'h66d3: y = 16'h200;
			16'h66d4: y = 16'h200;
			16'h66d5: y = 16'h200;
			16'h66d6: y = 16'h200;
			16'h66d7: y = 16'h200;
			16'h66d8: y = 16'h200;
			16'h66d9: y = 16'h200;
			16'h66da: y = 16'h200;
			16'h66db: y = 16'h200;
			16'h66dc: y = 16'h200;
			16'h66dd: y = 16'h200;
			16'h66de: y = 16'h200;
			16'h66df: y = 16'h200;
			16'h66e0: y = 16'h200;
			16'h66e1: y = 16'h200;
			16'h66e2: y = 16'h200;
			16'h66e3: y = 16'h200;
			16'h66e4: y = 16'h200;
			16'h66e5: y = 16'h200;
			16'h66e6: y = 16'h200;
			16'h66e7: y = 16'h200;
			16'h66e8: y = 16'h200;
			16'h66e9: y = 16'h200;
			16'h66ea: y = 16'h200;
			16'h66eb: y = 16'h200;
			16'h66ec: y = 16'h200;
			16'h66ed: y = 16'h200;
			16'h66ee: y = 16'h200;
			16'h66ef: y = 16'h200;
			16'h66f0: y = 16'h200;
			16'h66f1: y = 16'h200;
			16'h66f2: y = 16'h200;
			16'h66f3: y = 16'h200;
			16'h66f4: y = 16'h200;
			16'h66f5: y = 16'h200;
			16'h66f6: y = 16'h200;
			16'h66f7: y = 16'h200;
			16'h66f8: y = 16'h200;
			16'h66f9: y = 16'h200;
			16'h66fa: y = 16'h200;
			16'h66fb: y = 16'h200;
			16'h66fc: y = 16'h200;
			16'h66fd: y = 16'h200;
			16'h66fe: y = 16'h200;
			16'h66ff: y = 16'h200;
			16'h6700: y = 16'h200;
			16'h6701: y = 16'h200;
			16'h6702: y = 16'h200;
			16'h6703: y = 16'h200;
			16'h6704: y = 16'h200;
			16'h6705: y = 16'h200;
			16'h6706: y = 16'h200;
			16'h6707: y = 16'h200;
			16'h6708: y = 16'h200;
			16'h6709: y = 16'h200;
			16'h670a: y = 16'h200;
			16'h670b: y = 16'h200;
			16'h670c: y = 16'h200;
			16'h670d: y = 16'h200;
			16'h670e: y = 16'h200;
			16'h670f: y = 16'h200;
			16'h6710: y = 16'h200;
			16'h6711: y = 16'h200;
			16'h6712: y = 16'h200;
			16'h6713: y = 16'h200;
			16'h6714: y = 16'h200;
			16'h6715: y = 16'h200;
			16'h6716: y = 16'h200;
			16'h6717: y = 16'h200;
			16'h6718: y = 16'h200;
			16'h6719: y = 16'h200;
			16'h671a: y = 16'h200;
			16'h671b: y = 16'h200;
			16'h671c: y = 16'h200;
			16'h671d: y = 16'h200;
			16'h671e: y = 16'h200;
			16'h671f: y = 16'h200;
			16'h6720: y = 16'h200;
			16'h6721: y = 16'h200;
			16'h6722: y = 16'h200;
			16'h6723: y = 16'h200;
			16'h6724: y = 16'h200;
			16'h6725: y = 16'h200;
			16'h6726: y = 16'h200;
			16'h6727: y = 16'h200;
			16'h6728: y = 16'h200;
			16'h6729: y = 16'h200;
			16'h672a: y = 16'h200;
			16'h672b: y = 16'h200;
			16'h672c: y = 16'h200;
			16'h672d: y = 16'h200;
			16'h672e: y = 16'h200;
			16'h672f: y = 16'h200;
			16'h6730: y = 16'h200;
			16'h6731: y = 16'h200;
			16'h6732: y = 16'h200;
			16'h6733: y = 16'h200;
			16'h6734: y = 16'h200;
			16'h6735: y = 16'h200;
			16'h6736: y = 16'h200;
			16'h6737: y = 16'h200;
			16'h6738: y = 16'h200;
			16'h6739: y = 16'h200;
			16'h673a: y = 16'h200;
			16'h673b: y = 16'h200;
			16'h673c: y = 16'h200;
			16'h673d: y = 16'h200;
			16'h673e: y = 16'h200;
			16'h673f: y = 16'h200;
			16'h6740: y = 16'h200;
			16'h6741: y = 16'h200;
			16'h6742: y = 16'h200;
			16'h6743: y = 16'h200;
			16'h6744: y = 16'h200;
			16'h6745: y = 16'h200;
			16'h6746: y = 16'h200;
			16'h6747: y = 16'h200;
			16'h6748: y = 16'h200;
			16'h6749: y = 16'h200;
			16'h674a: y = 16'h200;
			16'h674b: y = 16'h200;
			16'h674c: y = 16'h200;
			16'h674d: y = 16'h200;
			16'h674e: y = 16'h200;
			16'h674f: y = 16'h200;
			16'h6750: y = 16'h200;
			16'h6751: y = 16'h200;
			16'h6752: y = 16'h200;
			16'h6753: y = 16'h200;
			16'h6754: y = 16'h200;
			16'h6755: y = 16'h200;
			16'h6756: y = 16'h200;
			16'h6757: y = 16'h200;
			16'h6758: y = 16'h200;
			16'h6759: y = 16'h200;
			16'h675a: y = 16'h200;
			16'h675b: y = 16'h200;
			16'h675c: y = 16'h200;
			16'h675d: y = 16'h200;
			16'h675e: y = 16'h200;
			16'h675f: y = 16'h200;
			16'h6760: y = 16'h200;
			16'h6761: y = 16'h200;
			16'h6762: y = 16'h200;
			16'h6763: y = 16'h200;
			16'h6764: y = 16'h200;
			16'h6765: y = 16'h200;
			16'h6766: y = 16'h200;
			16'h6767: y = 16'h200;
			16'h6768: y = 16'h200;
			16'h6769: y = 16'h200;
			16'h676a: y = 16'h200;
			16'h676b: y = 16'h200;
			16'h676c: y = 16'h200;
			16'h676d: y = 16'h200;
			16'h676e: y = 16'h200;
			16'h676f: y = 16'h200;
			16'h6770: y = 16'h200;
			16'h6771: y = 16'h200;
			16'h6772: y = 16'h200;
			16'h6773: y = 16'h200;
			16'h6774: y = 16'h200;
			16'h6775: y = 16'h200;
			16'h6776: y = 16'h200;
			16'h6777: y = 16'h200;
			16'h6778: y = 16'h200;
			16'h6779: y = 16'h200;
			16'h677a: y = 16'h200;
			16'h677b: y = 16'h200;
			16'h677c: y = 16'h200;
			16'h677d: y = 16'h200;
			16'h677e: y = 16'h200;
			16'h677f: y = 16'h200;
			16'h6780: y = 16'h200;
			16'h6781: y = 16'h200;
			16'h6782: y = 16'h200;
			16'h6783: y = 16'h200;
			16'h6784: y = 16'h200;
			16'h6785: y = 16'h200;
			16'h6786: y = 16'h200;
			16'h6787: y = 16'h200;
			16'h6788: y = 16'h200;
			16'h6789: y = 16'h200;
			16'h678a: y = 16'h200;
			16'h678b: y = 16'h200;
			16'h678c: y = 16'h200;
			16'h678d: y = 16'h200;
			16'h678e: y = 16'h200;
			16'h678f: y = 16'h200;
			16'h6790: y = 16'h200;
			16'h6791: y = 16'h200;
			16'h6792: y = 16'h200;
			16'h6793: y = 16'h200;
			16'h6794: y = 16'h200;
			16'h6795: y = 16'h200;
			16'h6796: y = 16'h200;
			16'h6797: y = 16'h200;
			16'h6798: y = 16'h200;
			16'h6799: y = 16'h200;
			16'h679a: y = 16'h200;
			16'h679b: y = 16'h200;
			16'h679c: y = 16'h200;
			16'h679d: y = 16'h200;
			16'h679e: y = 16'h200;
			16'h679f: y = 16'h200;
			16'h67a0: y = 16'h200;
			16'h67a1: y = 16'h200;
			16'h67a2: y = 16'h200;
			16'h67a3: y = 16'h200;
			16'h67a4: y = 16'h200;
			16'h67a5: y = 16'h200;
			16'h67a6: y = 16'h200;
			16'h67a7: y = 16'h200;
			16'h67a8: y = 16'h200;
			16'h67a9: y = 16'h200;
			16'h67aa: y = 16'h200;
			16'h67ab: y = 16'h200;
			16'h67ac: y = 16'h200;
			16'h67ad: y = 16'h200;
			16'h67ae: y = 16'h200;
			16'h67af: y = 16'h200;
			16'h67b0: y = 16'h200;
			16'h67b1: y = 16'h200;
			16'h67b2: y = 16'h200;
			16'h67b3: y = 16'h200;
			16'h67b4: y = 16'h200;
			16'h67b5: y = 16'h200;
			16'h67b6: y = 16'h200;
			16'h67b7: y = 16'h200;
			16'h67b8: y = 16'h200;
			16'h67b9: y = 16'h200;
			16'h67ba: y = 16'h200;
			16'h67bb: y = 16'h200;
			16'h67bc: y = 16'h200;
			16'h67bd: y = 16'h200;
			16'h67be: y = 16'h200;
			16'h67bf: y = 16'h200;
			16'h67c0: y = 16'h200;
			16'h67c1: y = 16'h200;
			16'h67c2: y = 16'h200;
			16'h67c3: y = 16'h200;
			16'h67c4: y = 16'h200;
			16'h67c5: y = 16'h200;
			16'h67c6: y = 16'h200;
			16'h67c7: y = 16'h200;
			16'h67c8: y = 16'h200;
			16'h67c9: y = 16'h200;
			16'h67ca: y = 16'h200;
			16'h67cb: y = 16'h200;
			16'h67cc: y = 16'h200;
			16'h67cd: y = 16'h200;
			16'h67ce: y = 16'h200;
			16'h67cf: y = 16'h200;
			16'h67d0: y = 16'h200;
			16'h67d1: y = 16'h200;
			16'h67d2: y = 16'h200;
			16'h67d3: y = 16'h200;
			16'h67d4: y = 16'h200;
			16'h67d5: y = 16'h200;
			16'h67d6: y = 16'h200;
			16'h67d7: y = 16'h200;
			16'h67d8: y = 16'h200;
			16'h67d9: y = 16'h200;
			16'h67da: y = 16'h200;
			16'h67db: y = 16'h200;
			16'h67dc: y = 16'h200;
			16'h67dd: y = 16'h200;
			16'h67de: y = 16'h200;
			16'h67df: y = 16'h200;
			16'h67e0: y = 16'h200;
			16'h67e1: y = 16'h200;
			16'h67e2: y = 16'h200;
			16'h67e3: y = 16'h200;
			16'h67e4: y = 16'h200;
			16'h67e5: y = 16'h200;
			16'h67e6: y = 16'h200;
			16'h67e7: y = 16'h200;
			16'h67e8: y = 16'h200;
			16'h67e9: y = 16'h200;
			16'h67ea: y = 16'h200;
			16'h67eb: y = 16'h200;
			16'h67ec: y = 16'h200;
			16'h67ed: y = 16'h200;
			16'h67ee: y = 16'h200;
			16'h67ef: y = 16'h200;
			16'h67f0: y = 16'h200;
			16'h67f1: y = 16'h200;
			16'h67f2: y = 16'h200;
			16'h67f3: y = 16'h200;
			16'h67f4: y = 16'h200;
			16'h67f5: y = 16'h200;
			16'h67f6: y = 16'h200;
			16'h67f7: y = 16'h200;
			16'h67f8: y = 16'h200;
			16'h67f9: y = 16'h200;
			16'h67fa: y = 16'h200;
			16'h67fb: y = 16'h200;
			16'h67fc: y = 16'h200;
			16'h67fd: y = 16'h200;
			16'h67fe: y = 16'h200;
			16'h67ff: y = 16'h200;
			16'h6800: y = 16'h200;
			16'h6801: y = 16'h200;
			16'h6802: y = 16'h200;
			16'h6803: y = 16'h200;
			16'h6804: y = 16'h200;
			16'h6805: y = 16'h200;
			16'h6806: y = 16'h200;
			16'h6807: y = 16'h200;
			16'h6808: y = 16'h200;
			16'h6809: y = 16'h200;
			16'h680a: y = 16'h200;
			16'h680b: y = 16'h200;
			16'h680c: y = 16'h200;
			16'h680d: y = 16'h200;
			16'h680e: y = 16'h200;
			16'h680f: y = 16'h200;
			16'h6810: y = 16'h200;
			16'h6811: y = 16'h200;
			16'h6812: y = 16'h200;
			16'h6813: y = 16'h200;
			16'h6814: y = 16'h200;
			16'h6815: y = 16'h200;
			16'h6816: y = 16'h200;
			16'h6817: y = 16'h200;
			16'h6818: y = 16'h200;
			16'h6819: y = 16'h200;
			16'h681a: y = 16'h200;
			16'h681b: y = 16'h200;
			16'h681c: y = 16'h200;
			16'h681d: y = 16'h200;
			16'h681e: y = 16'h200;
			16'h681f: y = 16'h200;
			16'h6820: y = 16'h200;
			16'h6821: y = 16'h200;
			16'h6822: y = 16'h200;
			16'h6823: y = 16'h200;
			16'h6824: y = 16'h200;
			16'h6825: y = 16'h200;
			16'h6826: y = 16'h200;
			16'h6827: y = 16'h200;
			16'h6828: y = 16'h200;
			16'h6829: y = 16'h200;
			16'h682a: y = 16'h200;
			16'h682b: y = 16'h200;
			16'h682c: y = 16'h200;
			16'h682d: y = 16'h200;
			16'h682e: y = 16'h200;
			16'h682f: y = 16'h200;
			16'h6830: y = 16'h200;
			16'h6831: y = 16'h200;
			16'h6832: y = 16'h200;
			16'h6833: y = 16'h200;
			16'h6834: y = 16'h200;
			16'h6835: y = 16'h200;
			16'h6836: y = 16'h200;
			16'h6837: y = 16'h200;
			16'h6838: y = 16'h200;
			16'h6839: y = 16'h200;
			16'h683a: y = 16'h200;
			16'h683b: y = 16'h200;
			16'h683c: y = 16'h200;
			16'h683d: y = 16'h200;
			16'h683e: y = 16'h200;
			16'h683f: y = 16'h200;
			16'h6840: y = 16'h200;
			16'h6841: y = 16'h200;
			16'h6842: y = 16'h200;
			16'h6843: y = 16'h200;
			16'h6844: y = 16'h200;
			16'h6845: y = 16'h200;
			16'h6846: y = 16'h200;
			16'h6847: y = 16'h200;
			16'h6848: y = 16'h200;
			16'h6849: y = 16'h200;
			16'h684a: y = 16'h200;
			16'h684b: y = 16'h200;
			16'h684c: y = 16'h200;
			16'h684d: y = 16'h200;
			16'h684e: y = 16'h200;
			16'h684f: y = 16'h200;
			16'h6850: y = 16'h200;
			16'h6851: y = 16'h200;
			16'h6852: y = 16'h200;
			16'h6853: y = 16'h200;
			16'h6854: y = 16'h200;
			16'h6855: y = 16'h200;
			16'h6856: y = 16'h200;
			16'h6857: y = 16'h200;
			16'h6858: y = 16'h200;
			16'h6859: y = 16'h200;
			16'h685a: y = 16'h200;
			16'h685b: y = 16'h200;
			16'h685c: y = 16'h200;
			16'h685d: y = 16'h200;
			16'h685e: y = 16'h200;
			16'h685f: y = 16'h200;
			16'h6860: y = 16'h200;
			16'h6861: y = 16'h200;
			16'h6862: y = 16'h200;
			16'h6863: y = 16'h200;
			16'h6864: y = 16'h200;
			16'h6865: y = 16'h200;
			16'h6866: y = 16'h200;
			16'h6867: y = 16'h200;
			16'h6868: y = 16'h200;
			16'h6869: y = 16'h200;
			16'h686a: y = 16'h200;
			16'h686b: y = 16'h200;
			16'h686c: y = 16'h200;
			16'h686d: y = 16'h200;
			16'h686e: y = 16'h200;
			16'h686f: y = 16'h200;
			16'h6870: y = 16'h200;
			16'h6871: y = 16'h200;
			16'h6872: y = 16'h200;
			16'h6873: y = 16'h200;
			16'h6874: y = 16'h200;
			16'h6875: y = 16'h200;
			16'h6876: y = 16'h200;
			16'h6877: y = 16'h200;
			16'h6878: y = 16'h200;
			16'h6879: y = 16'h200;
			16'h687a: y = 16'h200;
			16'h687b: y = 16'h200;
			16'h687c: y = 16'h200;
			16'h687d: y = 16'h200;
			16'h687e: y = 16'h200;
			16'h687f: y = 16'h200;
			16'h6880: y = 16'h200;
			16'h6881: y = 16'h200;
			16'h6882: y = 16'h200;
			16'h6883: y = 16'h200;
			16'h6884: y = 16'h200;
			16'h6885: y = 16'h200;
			16'h6886: y = 16'h200;
			16'h6887: y = 16'h200;
			16'h6888: y = 16'h200;
			16'h6889: y = 16'h200;
			16'h688a: y = 16'h200;
			16'h688b: y = 16'h200;
			16'h688c: y = 16'h200;
			16'h688d: y = 16'h200;
			16'h688e: y = 16'h200;
			16'h688f: y = 16'h200;
			16'h6890: y = 16'h200;
			16'h6891: y = 16'h200;
			16'h6892: y = 16'h200;
			16'h6893: y = 16'h200;
			16'h6894: y = 16'h200;
			16'h6895: y = 16'h200;
			16'h6896: y = 16'h200;
			16'h6897: y = 16'h200;
			16'h6898: y = 16'h200;
			16'h6899: y = 16'h200;
			16'h689a: y = 16'h200;
			16'h689b: y = 16'h200;
			16'h689c: y = 16'h200;
			16'h689d: y = 16'h200;
			16'h689e: y = 16'h200;
			16'h689f: y = 16'h200;
			16'h68a0: y = 16'h200;
			16'h68a1: y = 16'h200;
			16'h68a2: y = 16'h200;
			16'h68a3: y = 16'h200;
			16'h68a4: y = 16'h200;
			16'h68a5: y = 16'h200;
			16'h68a6: y = 16'h200;
			16'h68a7: y = 16'h200;
			16'h68a8: y = 16'h200;
			16'h68a9: y = 16'h200;
			16'h68aa: y = 16'h200;
			16'h68ab: y = 16'h200;
			16'h68ac: y = 16'h200;
			16'h68ad: y = 16'h200;
			16'h68ae: y = 16'h200;
			16'h68af: y = 16'h200;
			16'h68b0: y = 16'h200;
			16'h68b1: y = 16'h200;
			16'h68b2: y = 16'h200;
			16'h68b3: y = 16'h200;
			16'h68b4: y = 16'h200;
			16'h68b5: y = 16'h200;
			16'h68b6: y = 16'h200;
			16'h68b7: y = 16'h200;
			16'h68b8: y = 16'h200;
			16'h68b9: y = 16'h200;
			16'h68ba: y = 16'h200;
			16'h68bb: y = 16'h200;
			16'h68bc: y = 16'h200;
			16'h68bd: y = 16'h200;
			16'h68be: y = 16'h200;
			16'h68bf: y = 16'h200;
			16'h68c0: y = 16'h200;
			16'h68c1: y = 16'h200;
			16'h68c2: y = 16'h200;
			16'h68c3: y = 16'h200;
			16'h68c4: y = 16'h200;
			16'h68c5: y = 16'h200;
			16'h68c6: y = 16'h200;
			16'h68c7: y = 16'h200;
			16'h68c8: y = 16'h200;
			16'h68c9: y = 16'h200;
			16'h68ca: y = 16'h200;
			16'h68cb: y = 16'h200;
			16'h68cc: y = 16'h200;
			16'h68cd: y = 16'h200;
			16'h68ce: y = 16'h200;
			16'h68cf: y = 16'h200;
			16'h68d0: y = 16'h200;
			16'h68d1: y = 16'h200;
			16'h68d2: y = 16'h200;
			16'h68d3: y = 16'h200;
			16'h68d4: y = 16'h200;
			16'h68d5: y = 16'h200;
			16'h68d6: y = 16'h200;
			16'h68d7: y = 16'h200;
			16'h68d8: y = 16'h200;
			16'h68d9: y = 16'h200;
			16'h68da: y = 16'h200;
			16'h68db: y = 16'h200;
			16'h68dc: y = 16'h200;
			16'h68dd: y = 16'h200;
			16'h68de: y = 16'h200;
			16'h68df: y = 16'h200;
			16'h68e0: y = 16'h200;
			16'h68e1: y = 16'h200;
			16'h68e2: y = 16'h200;
			16'h68e3: y = 16'h200;
			16'h68e4: y = 16'h200;
			16'h68e5: y = 16'h200;
			16'h68e6: y = 16'h200;
			16'h68e7: y = 16'h200;
			16'h68e8: y = 16'h200;
			16'h68e9: y = 16'h200;
			16'h68ea: y = 16'h200;
			16'h68eb: y = 16'h200;
			16'h68ec: y = 16'h200;
			16'h68ed: y = 16'h200;
			16'h68ee: y = 16'h200;
			16'h68ef: y = 16'h200;
			16'h68f0: y = 16'h200;
			16'h68f1: y = 16'h200;
			16'h68f2: y = 16'h200;
			16'h68f3: y = 16'h200;
			16'h68f4: y = 16'h200;
			16'h68f5: y = 16'h200;
			16'h68f6: y = 16'h200;
			16'h68f7: y = 16'h200;
			16'h68f8: y = 16'h200;
			16'h68f9: y = 16'h200;
			16'h68fa: y = 16'h200;
			16'h68fb: y = 16'h200;
			16'h68fc: y = 16'h200;
			16'h68fd: y = 16'h200;
			16'h68fe: y = 16'h200;
			16'h68ff: y = 16'h200;
			16'h6900: y = 16'h200;
			16'h6901: y = 16'h200;
			16'h6902: y = 16'h200;
			16'h6903: y = 16'h200;
			16'h6904: y = 16'h200;
			16'h6905: y = 16'h200;
			16'h6906: y = 16'h200;
			16'h6907: y = 16'h200;
			16'h6908: y = 16'h200;
			16'h6909: y = 16'h200;
			16'h690a: y = 16'h200;
			16'h690b: y = 16'h200;
			16'h690c: y = 16'h200;
			16'h690d: y = 16'h200;
			16'h690e: y = 16'h200;
			16'h690f: y = 16'h200;
			16'h6910: y = 16'h200;
			16'h6911: y = 16'h200;
			16'h6912: y = 16'h200;
			16'h6913: y = 16'h200;
			16'h6914: y = 16'h200;
			16'h6915: y = 16'h200;
			16'h6916: y = 16'h200;
			16'h6917: y = 16'h200;
			16'h6918: y = 16'h200;
			16'h6919: y = 16'h200;
			16'h691a: y = 16'h200;
			16'h691b: y = 16'h200;
			16'h691c: y = 16'h200;
			16'h691d: y = 16'h200;
			16'h691e: y = 16'h200;
			16'h691f: y = 16'h200;
			16'h6920: y = 16'h200;
			16'h6921: y = 16'h200;
			16'h6922: y = 16'h200;
			16'h6923: y = 16'h200;
			16'h6924: y = 16'h200;
			16'h6925: y = 16'h200;
			16'h6926: y = 16'h200;
			16'h6927: y = 16'h200;
			16'h6928: y = 16'h200;
			16'h6929: y = 16'h200;
			16'h692a: y = 16'h200;
			16'h692b: y = 16'h200;
			16'h692c: y = 16'h200;
			16'h692d: y = 16'h200;
			16'h692e: y = 16'h200;
			16'h692f: y = 16'h200;
			16'h6930: y = 16'h200;
			16'h6931: y = 16'h200;
			16'h6932: y = 16'h200;
			16'h6933: y = 16'h200;
			16'h6934: y = 16'h200;
			16'h6935: y = 16'h200;
			16'h6936: y = 16'h200;
			16'h6937: y = 16'h200;
			16'h6938: y = 16'h200;
			16'h6939: y = 16'h200;
			16'h693a: y = 16'h200;
			16'h693b: y = 16'h200;
			16'h693c: y = 16'h200;
			16'h693d: y = 16'h200;
			16'h693e: y = 16'h200;
			16'h693f: y = 16'h200;
			16'h6940: y = 16'h200;
			16'h6941: y = 16'h200;
			16'h6942: y = 16'h200;
			16'h6943: y = 16'h200;
			16'h6944: y = 16'h200;
			16'h6945: y = 16'h200;
			16'h6946: y = 16'h200;
			16'h6947: y = 16'h200;
			16'h6948: y = 16'h200;
			16'h6949: y = 16'h200;
			16'h694a: y = 16'h200;
			16'h694b: y = 16'h200;
			16'h694c: y = 16'h200;
			16'h694d: y = 16'h200;
			16'h694e: y = 16'h200;
			16'h694f: y = 16'h200;
			16'h6950: y = 16'h200;
			16'h6951: y = 16'h200;
			16'h6952: y = 16'h200;
			16'h6953: y = 16'h200;
			16'h6954: y = 16'h200;
			16'h6955: y = 16'h200;
			16'h6956: y = 16'h200;
			16'h6957: y = 16'h200;
			16'h6958: y = 16'h200;
			16'h6959: y = 16'h200;
			16'h695a: y = 16'h200;
			16'h695b: y = 16'h200;
			16'h695c: y = 16'h200;
			16'h695d: y = 16'h200;
			16'h695e: y = 16'h200;
			16'h695f: y = 16'h200;
			16'h6960: y = 16'h200;
			16'h6961: y = 16'h200;
			16'h6962: y = 16'h200;
			16'h6963: y = 16'h200;
			16'h6964: y = 16'h200;
			16'h6965: y = 16'h200;
			16'h6966: y = 16'h200;
			16'h6967: y = 16'h200;
			16'h6968: y = 16'h200;
			16'h6969: y = 16'h200;
			16'h696a: y = 16'h200;
			16'h696b: y = 16'h200;
			16'h696c: y = 16'h200;
			16'h696d: y = 16'h200;
			16'h696e: y = 16'h200;
			16'h696f: y = 16'h200;
			16'h6970: y = 16'h200;
			16'h6971: y = 16'h200;
			16'h6972: y = 16'h200;
			16'h6973: y = 16'h200;
			16'h6974: y = 16'h200;
			16'h6975: y = 16'h200;
			16'h6976: y = 16'h200;
			16'h6977: y = 16'h200;
			16'h6978: y = 16'h200;
			16'h6979: y = 16'h200;
			16'h697a: y = 16'h200;
			16'h697b: y = 16'h200;
			16'h697c: y = 16'h200;
			16'h697d: y = 16'h200;
			16'h697e: y = 16'h200;
			16'h697f: y = 16'h200;
			16'h6980: y = 16'h200;
			16'h6981: y = 16'h200;
			16'h6982: y = 16'h200;
			16'h6983: y = 16'h200;
			16'h6984: y = 16'h200;
			16'h6985: y = 16'h200;
			16'h6986: y = 16'h200;
			16'h6987: y = 16'h200;
			16'h6988: y = 16'h200;
			16'h6989: y = 16'h200;
			16'h698a: y = 16'h200;
			16'h698b: y = 16'h200;
			16'h698c: y = 16'h200;
			16'h698d: y = 16'h200;
			16'h698e: y = 16'h200;
			16'h698f: y = 16'h200;
			16'h6990: y = 16'h200;
			16'h6991: y = 16'h200;
			16'h6992: y = 16'h200;
			16'h6993: y = 16'h200;
			16'h6994: y = 16'h200;
			16'h6995: y = 16'h200;
			16'h6996: y = 16'h200;
			16'h6997: y = 16'h200;
			16'h6998: y = 16'h200;
			16'h6999: y = 16'h200;
			16'h699a: y = 16'h200;
			16'h699b: y = 16'h200;
			16'h699c: y = 16'h200;
			16'h699d: y = 16'h200;
			16'h699e: y = 16'h200;
			16'h699f: y = 16'h200;
			16'h69a0: y = 16'h200;
			16'h69a1: y = 16'h200;
			16'h69a2: y = 16'h200;
			16'h69a3: y = 16'h200;
			16'h69a4: y = 16'h200;
			16'h69a5: y = 16'h200;
			16'h69a6: y = 16'h200;
			16'h69a7: y = 16'h200;
			16'h69a8: y = 16'h200;
			16'h69a9: y = 16'h200;
			16'h69aa: y = 16'h200;
			16'h69ab: y = 16'h200;
			16'h69ac: y = 16'h200;
			16'h69ad: y = 16'h200;
			16'h69ae: y = 16'h200;
			16'h69af: y = 16'h200;
			16'h69b0: y = 16'h200;
			16'h69b1: y = 16'h200;
			16'h69b2: y = 16'h200;
			16'h69b3: y = 16'h200;
			16'h69b4: y = 16'h200;
			16'h69b5: y = 16'h200;
			16'h69b6: y = 16'h200;
			16'h69b7: y = 16'h200;
			16'h69b8: y = 16'h200;
			16'h69b9: y = 16'h200;
			16'h69ba: y = 16'h200;
			16'h69bb: y = 16'h200;
			16'h69bc: y = 16'h200;
			16'h69bd: y = 16'h200;
			16'h69be: y = 16'h200;
			16'h69bf: y = 16'h200;
			16'h69c0: y = 16'h200;
			16'h69c1: y = 16'h200;
			16'h69c2: y = 16'h200;
			16'h69c3: y = 16'h200;
			16'h69c4: y = 16'h200;
			16'h69c5: y = 16'h200;
			16'h69c6: y = 16'h200;
			16'h69c7: y = 16'h200;
			16'h69c8: y = 16'h200;
			16'h69c9: y = 16'h200;
			16'h69ca: y = 16'h200;
			16'h69cb: y = 16'h200;
			16'h69cc: y = 16'h200;
			16'h69cd: y = 16'h200;
			16'h69ce: y = 16'h200;
			16'h69cf: y = 16'h200;
			16'h69d0: y = 16'h200;
			16'h69d1: y = 16'h200;
			16'h69d2: y = 16'h200;
			16'h69d3: y = 16'h200;
			16'h69d4: y = 16'h200;
			16'h69d5: y = 16'h200;
			16'h69d6: y = 16'h200;
			16'h69d7: y = 16'h200;
			16'h69d8: y = 16'h200;
			16'h69d9: y = 16'h200;
			16'h69da: y = 16'h200;
			16'h69db: y = 16'h200;
			16'h69dc: y = 16'h200;
			16'h69dd: y = 16'h200;
			16'h69de: y = 16'h200;
			16'h69df: y = 16'h200;
			16'h69e0: y = 16'h200;
			16'h69e1: y = 16'h200;
			16'h69e2: y = 16'h200;
			16'h69e3: y = 16'h200;
			16'h69e4: y = 16'h200;
			16'h69e5: y = 16'h200;
			16'h69e6: y = 16'h200;
			16'h69e7: y = 16'h200;
			16'h69e8: y = 16'h200;
			16'h69e9: y = 16'h200;
			16'h69ea: y = 16'h200;
			16'h69eb: y = 16'h200;
			16'h69ec: y = 16'h200;
			16'h69ed: y = 16'h200;
			16'h69ee: y = 16'h200;
			16'h69ef: y = 16'h200;
			16'h69f0: y = 16'h200;
			16'h69f1: y = 16'h200;
			16'h69f2: y = 16'h200;
			16'h69f3: y = 16'h200;
			16'h69f4: y = 16'h200;
			16'h69f5: y = 16'h200;
			16'h69f6: y = 16'h200;
			16'h69f7: y = 16'h200;
			16'h69f8: y = 16'h200;
			16'h69f9: y = 16'h200;
			16'h69fa: y = 16'h200;
			16'h69fb: y = 16'h200;
			16'h69fc: y = 16'h200;
			16'h69fd: y = 16'h200;
			16'h69fe: y = 16'h200;
			16'h69ff: y = 16'h200;
			16'h6a00: y = 16'h200;
			16'h6a01: y = 16'h200;
			16'h6a02: y = 16'h200;
			16'h6a03: y = 16'h200;
			16'h6a04: y = 16'h200;
			16'h6a05: y = 16'h200;
			16'h6a06: y = 16'h200;
			16'h6a07: y = 16'h200;
			16'h6a08: y = 16'h200;
			16'h6a09: y = 16'h200;
			16'h6a0a: y = 16'h200;
			16'h6a0b: y = 16'h200;
			16'h6a0c: y = 16'h200;
			16'h6a0d: y = 16'h200;
			16'h6a0e: y = 16'h200;
			16'h6a0f: y = 16'h200;
			16'h6a10: y = 16'h200;
			16'h6a11: y = 16'h200;
			16'h6a12: y = 16'h200;
			16'h6a13: y = 16'h200;
			16'h6a14: y = 16'h200;
			16'h6a15: y = 16'h200;
			16'h6a16: y = 16'h200;
			16'h6a17: y = 16'h200;
			16'h6a18: y = 16'h200;
			16'h6a19: y = 16'h200;
			16'h6a1a: y = 16'h200;
			16'h6a1b: y = 16'h200;
			16'h6a1c: y = 16'h200;
			16'h6a1d: y = 16'h200;
			16'h6a1e: y = 16'h200;
			16'h6a1f: y = 16'h200;
			16'h6a20: y = 16'h200;
			16'h6a21: y = 16'h200;
			16'h6a22: y = 16'h200;
			16'h6a23: y = 16'h200;
			16'h6a24: y = 16'h200;
			16'h6a25: y = 16'h200;
			16'h6a26: y = 16'h200;
			16'h6a27: y = 16'h200;
			16'h6a28: y = 16'h200;
			16'h6a29: y = 16'h200;
			16'h6a2a: y = 16'h200;
			16'h6a2b: y = 16'h200;
			16'h6a2c: y = 16'h200;
			16'h6a2d: y = 16'h200;
			16'h6a2e: y = 16'h200;
			16'h6a2f: y = 16'h200;
			16'h6a30: y = 16'h200;
			16'h6a31: y = 16'h200;
			16'h6a32: y = 16'h200;
			16'h6a33: y = 16'h200;
			16'h6a34: y = 16'h200;
			16'h6a35: y = 16'h200;
			16'h6a36: y = 16'h200;
			16'h6a37: y = 16'h200;
			16'h6a38: y = 16'h200;
			16'h6a39: y = 16'h200;
			16'h6a3a: y = 16'h200;
			16'h6a3b: y = 16'h200;
			16'h6a3c: y = 16'h200;
			16'h6a3d: y = 16'h200;
			16'h6a3e: y = 16'h200;
			16'h6a3f: y = 16'h200;
			16'h6a40: y = 16'h200;
			16'h6a41: y = 16'h200;
			16'h6a42: y = 16'h200;
			16'h6a43: y = 16'h200;
			16'h6a44: y = 16'h200;
			16'h6a45: y = 16'h200;
			16'h6a46: y = 16'h200;
			16'h6a47: y = 16'h200;
			16'h6a48: y = 16'h200;
			16'h6a49: y = 16'h200;
			16'h6a4a: y = 16'h200;
			16'h6a4b: y = 16'h200;
			16'h6a4c: y = 16'h200;
			16'h6a4d: y = 16'h200;
			16'h6a4e: y = 16'h200;
			16'h6a4f: y = 16'h200;
			16'h6a50: y = 16'h200;
			16'h6a51: y = 16'h200;
			16'h6a52: y = 16'h200;
			16'h6a53: y = 16'h200;
			16'h6a54: y = 16'h200;
			16'h6a55: y = 16'h200;
			16'h6a56: y = 16'h200;
			16'h6a57: y = 16'h200;
			16'h6a58: y = 16'h200;
			16'h6a59: y = 16'h200;
			16'h6a5a: y = 16'h200;
			16'h6a5b: y = 16'h200;
			16'h6a5c: y = 16'h200;
			16'h6a5d: y = 16'h200;
			16'h6a5e: y = 16'h200;
			16'h6a5f: y = 16'h200;
			16'h6a60: y = 16'h200;
			16'h6a61: y = 16'h200;
			16'h6a62: y = 16'h200;
			16'h6a63: y = 16'h200;
			16'h6a64: y = 16'h200;
			16'h6a65: y = 16'h200;
			16'h6a66: y = 16'h200;
			16'h6a67: y = 16'h200;
			16'h6a68: y = 16'h200;
			16'h6a69: y = 16'h200;
			16'h6a6a: y = 16'h200;
			16'h6a6b: y = 16'h200;
			16'h6a6c: y = 16'h200;
			16'h6a6d: y = 16'h200;
			16'h6a6e: y = 16'h200;
			16'h6a6f: y = 16'h200;
			16'h6a70: y = 16'h200;
			16'h6a71: y = 16'h200;
			16'h6a72: y = 16'h200;
			16'h6a73: y = 16'h200;
			16'h6a74: y = 16'h200;
			16'h6a75: y = 16'h200;
			16'h6a76: y = 16'h200;
			16'h6a77: y = 16'h200;
			16'h6a78: y = 16'h200;
			16'h6a79: y = 16'h200;
			16'h6a7a: y = 16'h200;
			16'h6a7b: y = 16'h200;
			16'h6a7c: y = 16'h200;
			16'h6a7d: y = 16'h200;
			16'h6a7e: y = 16'h200;
			16'h6a7f: y = 16'h200;
			16'h6a80: y = 16'h200;
			16'h6a81: y = 16'h200;
			16'h6a82: y = 16'h200;
			16'h6a83: y = 16'h200;
			16'h6a84: y = 16'h200;
			16'h6a85: y = 16'h200;
			16'h6a86: y = 16'h200;
			16'h6a87: y = 16'h200;
			16'h6a88: y = 16'h200;
			16'h6a89: y = 16'h200;
			16'h6a8a: y = 16'h200;
			16'h6a8b: y = 16'h200;
			16'h6a8c: y = 16'h200;
			16'h6a8d: y = 16'h200;
			16'h6a8e: y = 16'h200;
			16'h6a8f: y = 16'h200;
			16'h6a90: y = 16'h200;
			16'h6a91: y = 16'h200;
			16'h6a92: y = 16'h200;
			16'h6a93: y = 16'h200;
			16'h6a94: y = 16'h200;
			16'h6a95: y = 16'h200;
			16'h6a96: y = 16'h200;
			16'h6a97: y = 16'h200;
			16'h6a98: y = 16'h200;
			16'h6a99: y = 16'h200;
			16'h6a9a: y = 16'h200;
			16'h6a9b: y = 16'h200;
			16'h6a9c: y = 16'h200;
			16'h6a9d: y = 16'h200;
			16'h6a9e: y = 16'h200;
			16'h6a9f: y = 16'h200;
			16'h6aa0: y = 16'h200;
			16'h6aa1: y = 16'h200;
			16'h6aa2: y = 16'h200;
			16'h6aa3: y = 16'h200;
			16'h6aa4: y = 16'h200;
			16'h6aa5: y = 16'h200;
			16'h6aa6: y = 16'h200;
			16'h6aa7: y = 16'h200;
			16'h6aa8: y = 16'h200;
			16'h6aa9: y = 16'h200;
			16'h6aaa: y = 16'h200;
			16'h6aab: y = 16'h200;
			16'h6aac: y = 16'h200;
			16'h6aad: y = 16'h200;
			16'h6aae: y = 16'h200;
			16'h6aaf: y = 16'h200;
			16'h6ab0: y = 16'h200;
			16'h6ab1: y = 16'h200;
			16'h6ab2: y = 16'h200;
			16'h6ab3: y = 16'h200;
			16'h6ab4: y = 16'h200;
			16'h6ab5: y = 16'h200;
			16'h6ab6: y = 16'h200;
			16'h6ab7: y = 16'h200;
			16'h6ab8: y = 16'h200;
			16'h6ab9: y = 16'h200;
			16'h6aba: y = 16'h200;
			16'h6abb: y = 16'h200;
			16'h6abc: y = 16'h200;
			16'h6abd: y = 16'h200;
			16'h6abe: y = 16'h200;
			16'h6abf: y = 16'h200;
			16'h6ac0: y = 16'h200;
			16'h6ac1: y = 16'h200;
			16'h6ac2: y = 16'h200;
			16'h6ac3: y = 16'h200;
			16'h6ac4: y = 16'h200;
			16'h6ac5: y = 16'h200;
			16'h6ac6: y = 16'h200;
			16'h6ac7: y = 16'h200;
			16'h6ac8: y = 16'h200;
			16'h6ac9: y = 16'h200;
			16'h6aca: y = 16'h200;
			16'h6acb: y = 16'h200;
			16'h6acc: y = 16'h200;
			16'h6acd: y = 16'h200;
			16'h6ace: y = 16'h200;
			16'h6acf: y = 16'h200;
			16'h6ad0: y = 16'h200;
			16'h6ad1: y = 16'h200;
			16'h6ad2: y = 16'h200;
			16'h6ad3: y = 16'h200;
			16'h6ad4: y = 16'h200;
			16'h6ad5: y = 16'h200;
			16'h6ad6: y = 16'h200;
			16'h6ad7: y = 16'h200;
			16'h6ad8: y = 16'h200;
			16'h6ad9: y = 16'h200;
			16'h6ada: y = 16'h200;
			16'h6adb: y = 16'h200;
			16'h6adc: y = 16'h200;
			16'h6add: y = 16'h200;
			16'h6ade: y = 16'h200;
			16'h6adf: y = 16'h200;
			16'h6ae0: y = 16'h200;
			16'h6ae1: y = 16'h200;
			16'h6ae2: y = 16'h200;
			16'h6ae3: y = 16'h200;
			16'h6ae4: y = 16'h200;
			16'h6ae5: y = 16'h200;
			16'h6ae6: y = 16'h200;
			16'h6ae7: y = 16'h200;
			16'h6ae8: y = 16'h200;
			16'h6ae9: y = 16'h200;
			16'h6aea: y = 16'h200;
			16'h6aeb: y = 16'h200;
			16'h6aec: y = 16'h200;
			16'h6aed: y = 16'h200;
			16'h6aee: y = 16'h200;
			16'h6aef: y = 16'h200;
			16'h6af0: y = 16'h200;
			16'h6af1: y = 16'h200;
			16'h6af2: y = 16'h200;
			16'h6af3: y = 16'h200;
			16'h6af4: y = 16'h200;
			16'h6af5: y = 16'h200;
			16'h6af6: y = 16'h200;
			16'h6af7: y = 16'h200;
			16'h6af8: y = 16'h200;
			16'h6af9: y = 16'h200;
			16'h6afa: y = 16'h200;
			16'h6afb: y = 16'h200;
			16'h6afc: y = 16'h200;
			16'h6afd: y = 16'h200;
			16'h6afe: y = 16'h200;
			16'h6aff: y = 16'h200;
			16'h6b00: y = 16'h200;
			16'h6b01: y = 16'h200;
			16'h6b02: y = 16'h200;
			16'h6b03: y = 16'h200;
			16'h6b04: y = 16'h200;
			16'h6b05: y = 16'h200;
			16'h6b06: y = 16'h200;
			16'h6b07: y = 16'h200;
			16'h6b08: y = 16'h200;
			16'h6b09: y = 16'h200;
			16'h6b0a: y = 16'h200;
			16'h6b0b: y = 16'h200;
			16'h6b0c: y = 16'h200;
			16'h6b0d: y = 16'h200;
			16'h6b0e: y = 16'h200;
			16'h6b0f: y = 16'h200;
			16'h6b10: y = 16'h200;
			16'h6b11: y = 16'h200;
			16'h6b12: y = 16'h200;
			16'h6b13: y = 16'h200;
			16'h6b14: y = 16'h200;
			16'h6b15: y = 16'h200;
			16'h6b16: y = 16'h200;
			16'h6b17: y = 16'h200;
			16'h6b18: y = 16'h200;
			16'h6b19: y = 16'h200;
			16'h6b1a: y = 16'h200;
			16'h6b1b: y = 16'h200;
			16'h6b1c: y = 16'h200;
			16'h6b1d: y = 16'h200;
			16'h6b1e: y = 16'h200;
			16'h6b1f: y = 16'h200;
			16'h6b20: y = 16'h200;
			16'h6b21: y = 16'h200;
			16'h6b22: y = 16'h200;
			16'h6b23: y = 16'h200;
			16'h6b24: y = 16'h200;
			16'h6b25: y = 16'h200;
			16'h6b26: y = 16'h200;
			16'h6b27: y = 16'h200;
			16'h6b28: y = 16'h200;
			16'h6b29: y = 16'h200;
			16'h6b2a: y = 16'h200;
			16'h6b2b: y = 16'h200;
			16'h6b2c: y = 16'h200;
			16'h6b2d: y = 16'h200;
			16'h6b2e: y = 16'h200;
			16'h6b2f: y = 16'h200;
			16'h6b30: y = 16'h200;
			16'h6b31: y = 16'h200;
			16'h6b32: y = 16'h200;
			16'h6b33: y = 16'h200;
			16'h6b34: y = 16'h200;
			16'h6b35: y = 16'h200;
			16'h6b36: y = 16'h200;
			16'h6b37: y = 16'h200;
			16'h6b38: y = 16'h200;
			16'h6b39: y = 16'h200;
			16'h6b3a: y = 16'h200;
			16'h6b3b: y = 16'h200;
			16'h6b3c: y = 16'h200;
			16'h6b3d: y = 16'h200;
			16'h6b3e: y = 16'h200;
			16'h6b3f: y = 16'h200;
			16'h6b40: y = 16'h200;
			16'h6b41: y = 16'h200;
			16'h6b42: y = 16'h200;
			16'h6b43: y = 16'h200;
			16'h6b44: y = 16'h200;
			16'h6b45: y = 16'h200;
			16'h6b46: y = 16'h200;
			16'h6b47: y = 16'h200;
			16'h6b48: y = 16'h200;
			16'h6b49: y = 16'h200;
			16'h6b4a: y = 16'h200;
			16'h6b4b: y = 16'h200;
			16'h6b4c: y = 16'h200;
			16'h6b4d: y = 16'h200;
			16'h6b4e: y = 16'h200;
			16'h6b4f: y = 16'h200;
			16'h6b50: y = 16'h200;
			16'h6b51: y = 16'h200;
			16'h6b52: y = 16'h200;
			16'h6b53: y = 16'h200;
			16'h6b54: y = 16'h200;
			16'h6b55: y = 16'h200;
			16'h6b56: y = 16'h200;
			16'h6b57: y = 16'h200;
			16'h6b58: y = 16'h200;
			16'h6b59: y = 16'h200;
			16'h6b5a: y = 16'h200;
			16'h6b5b: y = 16'h200;
			16'h6b5c: y = 16'h200;
			16'h6b5d: y = 16'h200;
			16'h6b5e: y = 16'h200;
			16'h6b5f: y = 16'h200;
			16'h6b60: y = 16'h200;
			16'h6b61: y = 16'h200;
			16'h6b62: y = 16'h200;
			16'h6b63: y = 16'h200;
			16'h6b64: y = 16'h200;
			16'h6b65: y = 16'h200;
			16'h6b66: y = 16'h200;
			16'h6b67: y = 16'h200;
			16'h6b68: y = 16'h200;
			16'h6b69: y = 16'h200;
			16'h6b6a: y = 16'h200;
			16'h6b6b: y = 16'h200;
			16'h6b6c: y = 16'h200;
			16'h6b6d: y = 16'h200;
			16'h6b6e: y = 16'h200;
			16'h6b6f: y = 16'h200;
			16'h6b70: y = 16'h200;
			16'h6b71: y = 16'h200;
			16'h6b72: y = 16'h200;
			16'h6b73: y = 16'h200;
			16'h6b74: y = 16'h200;
			16'h6b75: y = 16'h200;
			16'h6b76: y = 16'h200;
			16'h6b77: y = 16'h200;
			16'h6b78: y = 16'h200;
			16'h6b79: y = 16'h200;
			16'h6b7a: y = 16'h200;
			16'h6b7b: y = 16'h200;
			16'h6b7c: y = 16'h200;
			16'h6b7d: y = 16'h200;
			16'h6b7e: y = 16'h200;
			16'h6b7f: y = 16'h200;
			16'h6b80: y = 16'h200;
			16'h6b81: y = 16'h200;
			16'h6b82: y = 16'h200;
			16'h6b83: y = 16'h200;
			16'h6b84: y = 16'h200;
			16'h6b85: y = 16'h200;
			16'h6b86: y = 16'h200;
			16'h6b87: y = 16'h200;
			16'h6b88: y = 16'h200;
			16'h6b89: y = 16'h200;
			16'h6b8a: y = 16'h200;
			16'h6b8b: y = 16'h200;
			16'h6b8c: y = 16'h200;
			16'h6b8d: y = 16'h200;
			16'h6b8e: y = 16'h200;
			16'h6b8f: y = 16'h200;
			16'h6b90: y = 16'h200;
			16'h6b91: y = 16'h200;
			16'h6b92: y = 16'h200;
			16'h6b93: y = 16'h200;
			16'h6b94: y = 16'h200;
			16'h6b95: y = 16'h200;
			16'h6b96: y = 16'h200;
			16'h6b97: y = 16'h200;
			16'h6b98: y = 16'h200;
			16'h6b99: y = 16'h200;
			16'h6b9a: y = 16'h200;
			16'h6b9b: y = 16'h200;
			16'h6b9c: y = 16'h200;
			16'h6b9d: y = 16'h200;
			16'h6b9e: y = 16'h200;
			16'h6b9f: y = 16'h200;
			16'h6ba0: y = 16'h200;
			16'h6ba1: y = 16'h200;
			16'h6ba2: y = 16'h200;
			16'h6ba3: y = 16'h200;
			16'h6ba4: y = 16'h200;
			16'h6ba5: y = 16'h200;
			16'h6ba6: y = 16'h200;
			16'h6ba7: y = 16'h200;
			16'h6ba8: y = 16'h200;
			16'h6ba9: y = 16'h200;
			16'h6baa: y = 16'h200;
			16'h6bab: y = 16'h200;
			16'h6bac: y = 16'h200;
			16'h6bad: y = 16'h200;
			16'h6bae: y = 16'h200;
			16'h6baf: y = 16'h200;
			16'h6bb0: y = 16'h200;
			16'h6bb1: y = 16'h200;
			16'h6bb2: y = 16'h200;
			16'h6bb3: y = 16'h200;
			16'h6bb4: y = 16'h200;
			16'h6bb5: y = 16'h200;
			16'h6bb6: y = 16'h200;
			16'h6bb7: y = 16'h200;
			16'h6bb8: y = 16'h200;
			16'h6bb9: y = 16'h200;
			16'h6bba: y = 16'h200;
			16'h6bbb: y = 16'h200;
			16'h6bbc: y = 16'h200;
			16'h6bbd: y = 16'h200;
			16'h6bbe: y = 16'h200;
			16'h6bbf: y = 16'h200;
			16'h6bc0: y = 16'h200;
			16'h6bc1: y = 16'h200;
			16'h6bc2: y = 16'h200;
			16'h6bc3: y = 16'h200;
			16'h6bc4: y = 16'h200;
			16'h6bc5: y = 16'h200;
			16'h6bc6: y = 16'h200;
			16'h6bc7: y = 16'h200;
			16'h6bc8: y = 16'h200;
			16'h6bc9: y = 16'h200;
			16'h6bca: y = 16'h200;
			16'h6bcb: y = 16'h200;
			16'h6bcc: y = 16'h200;
			16'h6bcd: y = 16'h200;
			16'h6bce: y = 16'h200;
			16'h6bcf: y = 16'h200;
			16'h6bd0: y = 16'h200;
			16'h6bd1: y = 16'h200;
			16'h6bd2: y = 16'h200;
			16'h6bd3: y = 16'h200;
			16'h6bd4: y = 16'h200;
			16'h6bd5: y = 16'h200;
			16'h6bd6: y = 16'h200;
			16'h6bd7: y = 16'h200;
			16'h6bd8: y = 16'h200;
			16'h6bd9: y = 16'h200;
			16'h6bda: y = 16'h200;
			16'h6bdb: y = 16'h200;
			16'h6bdc: y = 16'h200;
			16'h6bdd: y = 16'h200;
			16'h6bde: y = 16'h200;
			16'h6bdf: y = 16'h200;
			16'h6be0: y = 16'h200;
			16'h6be1: y = 16'h200;
			16'h6be2: y = 16'h200;
			16'h6be3: y = 16'h200;
			16'h6be4: y = 16'h200;
			16'h6be5: y = 16'h200;
			16'h6be6: y = 16'h200;
			16'h6be7: y = 16'h200;
			16'h6be8: y = 16'h200;
			16'h6be9: y = 16'h200;
			16'h6bea: y = 16'h200;
			16'h6beb: y = 16'h200;
			16'h6bec: y = 16'h200;
			16'h6bed: y = 16'h200;
			16'h6bee: y = 16'h200;
			16'h6bef: y = 16'h200;
			16'h6bf0: y = 16'h200;
			16'h6bf1: y = 16'h200;
			16'h6bf2: y = 16'h200;
			16'h6bf3: y = 16'h200;
			16'h6bf4: y = 16'h200;
			16'h6bf5: y = 16'h200;
			16'h6bf6: y = 16'h200;
			16'h6bf7: y = 16'h200;
			16'h6bf8: y = 16'h200;
			16'h6bf9: y = 16'h200;
			16'h6bfa: y = 16'h200;
			16'h6bfb: y = 16'h200;
			16'h6bfc: y = 16'h200;
			16'h6bfd: y = 16'h200;
			16'h6bfe: y = 16'h200;
			16'h6bff: y = 16'h200;
			16'h6c00: y = 16'h200;
			16'h6c01: y = 16'h200;
			16'h6c02: y = 16'h200;
			16'h6c03: y = 16'h200;
			16'h6c04: y = 16'h200;
			16'h6c05: y = 16'h200;
			16'h6c06: y = 16'h200;
			16'h6c07: y = 16'h200;
			16'h6c08: y = 16'h200;
			16'h6c09: y = 16'h200;
			16'h6c0a: y = 16'h200;
			16'h6c0b: y = 16'h200;
			16'h6c0c: y = 16'h200;
			16'h6c0d: y = 16'h200;
			16'h6c0e: y = 16'h200;
			16'h6c0f: y = 16'h200;
			16'h6c10: y = 16'h200;
			16'h6c11: y = 16'h200;
			16'h6c12: y = 16'h200;
			16'h6c13: y = 16'h200;
			16'h6c14: y = 16'h200;
			16'h6c15: y = 16'h200;
			16'h6c16: y = 16'h200;
			16'h6c17: y = 16'h200;
			16'h6c18: y = 16'h200;
			16'h6c19: y = 16'h200;
			16'h6c1a: y = 16'h200;
			16'h6c1b: y = 16'h200;
			16'h6c1c: y = 16'h200;
			16'h6c1d: y = 16'h200;
			16'h6c1e: y = 16'h200;
			16'h6c1f: y = 16'h200;
			16'h6c20: y = 16'h200;
			16'h6c21: y = 16'h200;
			16'h6c22: y = 16'h200;
			16'h6c23: y = 16'h200;
			16'h6c24: y = 16'h200;
			16'h6c25: y = 16'h200;
			16'h6c26: y = 16'h200;
			16'h6c27: y = 16'h200;
			16'h6c28: y = 16'h200;
			16'h6c29: y = 16'h200;
			16'h6c2a: y = 16'h200;
			16'h6c2b: y = 16'h200;
			16'h6c2c: y = 16'h200;
			16'h6c2d: y = 16'h200;
			16'h6c2e: y = 16'h200;
			16'h6c2f: y = 16'h200;
			16'h6c30: y = 16'h200;
			16'h6c31: y = 16'h200;
			16'h6c32: y = 16'h200;
			16'h6c33: y = 16'h200;
			16'h6c34: y = 16'h200;
			16'h6c35: y = 16'h200;
			16'h6c36: y = 16'h200;
			16'h6c37: y = 16'h200;
			16'h6c38: y = 16'h200;
			16'h6c39: y = 16'h200;
			16'h6c3a: y = 16'h200;
			16'h6c3b: y = 16'h200;
			16'h6c3c: y = 16'h200;
			16'h6c3d: y = 16'h200;
			16'h6c3e: y = 16'h200;
			16'h6c3f: y = 16'h200;
			16'h6c40: y = 16'h200;
			16'h6c41: y = 16'h200;
			16'h6c42: y = 16'h200;
			16'h6c43: y = 16'h200;
			16'h6c44: y = 16'h200;
			16'h6c45: y = 16'h200;
			16'h6c46: y = 16'h200;
			16'h6c47: y = 16'h200;
			16'h6c48: y = 16'h200;
			16'h6c49: y = 16'h200;
			16'h6c4a: y = 16'h200;
			16'h6c4b: y = 16'h200;
			16'h6c4c: y = 16'h200;
			16'h6c4d: y = 16'h200;
			16'h6c4e: y = 16'h200;
			16'h6c4f: y = 16'h200;
			16'h6c50: y = 16'h200;
			16'h6c51: y = 16'h200;
			16'h6c52: y = 16'h200;
			16'h6c53: y = 16'h200;
			16'h6c54: y = 16'h200;
			16'h6c55: y = 16'h200;
			16'h6c56: y = 16'h200;
			16'h6c57: y = 16'h200;
			16'h6c58: y = 16'h200;
			16'h6c59: y = 16'h200;
			16'h6c5a: y = 16'h200;
			16'h6c5b: y = 16'h200;
			16'h6c5c: y = 16'h200;
			16'h6c5d: y = 16'h200;
			16'h6c5e: y = 16'h200;
			16'h6c5f: y = 16'h200;
			16'h6c60: y = 16'h200;
			16'h6c61: y = 16'h200;
			16'h6c62: y = 16'h200;
			16'h6c63: y = 16'h200;
			16'h6c64: y = 16'h200;
			16'h6c65: y = 16'h200;
			16'h6c66: y = 16'h200;
			16'h6c67: y = 16'h200;
			16'h6c68: y = 16'h200;
			16'h6c69: y = 16'h200;
			16'h6c6a: y = 16'h200;
			16'h6c6b: y = 16'h200;
			16'h6c6c: y = 16'h200;
			16'h6c6d: y = 16'h200;
			16'h6c6e: y = 16'h200;
			16'h6c6f: y = 16'h200;
			16'h6c70: y = 16'h200;
			16'h6c71: y = 16'h200;
			16'h6c72: y = 16'h200;
			16'h6c73: y = 16'h200;
			16'h6c74: y = 16'h200;
			16'h6c75: y = 16'h200;
			16'h6c76: y = 16'h200;
			16'h6c77: y = 16'h200;
			16'h6c78: y = 16'h200;
			16'h6c79: y = 16'h200;
			16'h6c7a: y = 16'h200;
			16'h6c7b: y = 16'h200;
			16'h6c7c: y = 16'h200;
			16'h6c7d: y = 16'h200;
			16'h6c7e: y = 16'h200;
			16'h6c7f: y = 16'h200;
			16'h6c80: y = 16'h200;
			16'h6c81: y = 16'h200;
			16'h6c82: y = 16'h200;
			16'h6c83: y = 16'h200;
			16'h6c84: y = 16'h200;
			16'h6c85: y = 16'h200;
			16'h6c86: y = 16'h200;
			16'h6c87: y = 16'h200;
			16'h6c88: y = 16'h200;
			16'h6c89: y = 16'h200;
			16'h6c8a: y = 16'h200;
			16'h6c8b: y = 16'h200;
			16'h6c8c: y = 16'h200;
			16'h6c8d: y = 16'h200;
			16'h6c8e: y = 16'h200;
			16'h6c8f: y = 16'h200;
			16'h6c90: y = 16'h200;
			16'h6c91: y = 16'h200;
			16'h6c92: y = 16'h200;
			16'h6c93: y = 16'h200;
			16'h6c94: y = 16'h200;
			16'h6c95: y = 16'h200;
			16'h6c96: y = 16'h200;
			16'h6c97: y = 16'h200;
			16'h6c98: y = 16'h200;
			16'h6c99: y = 16'h200;
			16'h6c9a: y = 16'h200;
			16'h6c9b: y = 16'h200;
			16'h6c9c: y = 16'h200;
			16'h6c9d: y = 16'h200;
			16'h6c9e: y = 16'h200;
			16'h6c9f: y = 16'h200;
			16'h6ca0: y = 16'h200;
			16'h6ca1: y = 16'h200;
			16'h6ca2: y = 16'h200;
			16'h6ca3: y = 16'h200;
			16'h6ca4: y = 16'h200;
			16'h6ca5: y = 16'h200;
			16'h6ca6: y = 16'h200;
			16'h6ca7: y = 16'h200;
			16'h6ca8: y = 16'h200;
			16'h6ca9: y = 16'h200;
			16'h6caa: y = 16'h200;
			16'h6cab: y = 16'h200;
			16'h6cac: y = 16'h200;
			16'h6cad: y = 16'h200;
			16'h6cae: y = 16'h200;
			16'h6caf: y = 16'h200;
			16'h6cb0: y = 16'h200;
			16'h6cb1: y = 16'h200;
			16'h6cb2: y = 16'h200;
			16'h6cb3: y = 16'h200;
			16'h6cb4: y = 16'h200;
			16'h6cb5: y = 16'h200;
			16'h6cb6: y = 16'h200;
			16'h6cb7: y = 16'h200;
			16'h6cb8: y = 16'h200;
			16'h6cb9: y = 16'h200;
			16'h6cba: y = 16'h200;
			16'h6cbb: y = 16'h200;
			16'h6cbc: y = 16'h200;
			16'h6cbd: y = 16'h200;
			16'h6cbe: y = 16'h200;
			16'h6cbf: y = 16'h200;
			16'h6cc0: y = 16'h200;
			16'h6cc1: y = 16'h200;
			16'h6cc2: y = 16'h200;
			16'h6cc3: y = 16'h200;
			16'h6cc4: y = 16'h200;
			16'h6cc5: y = 16'h200;
			16'h6cc6: y = 16'h200;
			16'h6cc7: y = 16'h200;
			16'h6cc8: y = 16'h200;
			16'h6cc9: y = 16'h200;
			16'h6cca: y = 16'h200;
			16'h6ccb: y = 16'h200;
			16'h6ccc: y = 16'h200;
			16'h6ccd: y = 16'h200;
			16'h6cce: y = 16'h200;
			16'h6ccf: y = 16'h200;
			16'h6cd0: y = 16'h200;
			16'h6cd1: y = 16'h200;
			16'h6cd2: y = 16'h200;
			16'h6cd3: y = 16'h200;
			16'h6cd4: y = 16'h200;
			16'h6cd5: y = 16'h200;
			16'h6cd6: y = 16'h200;
			16'h6cd7: y = 16'h200;
			16'h6cd8: y = 16'h200;
			16'h6cd9: y = 16'h200;
			16'h6cda: y = 16'h200;
			16'h6cdb: y = 16'h200;
			16'h6cdc: y = 16'h200;
			16'h6cdd: y = 16'h200;
			16'h6cde: y = 16'h200;
			16'h6cdf: y = 16'h200;
			16'h6ce0: y = 16'h200;
			16'h6ce1: y = 16'h200;
			16'h6ce2: y = 16'h200;
			16'h6ce3: y = 16'h200;
			16'h6ce4: y = 16'h200;
			16'h6ce5: y = 16'h200;
			16'h6ce6: y = 16'h200;
			16'h6ce7: y = 16'h200;
			16'h6ce8: y = 16'h200;
			16'h6ce9: y = 16'h200;
			16'h6cea: y = 16'h200;
			16'h6ceb: y = 16'h200;
			16'h6cec: y = 16'h200;
			16'h6ced: y = 16'h200;
			16'h6cee: y = 16'h200;
			16'h6cef: y = 16'h200;
			16'h6cf0: y = 16'h200;
			16'h6cf1: y = 16'h200;
			16'h6cf2: y = 16'h200;
			16'h6cf3: y = 16'h200;
			16'h6cf4: y = 16'h200;
			16'h6cf5: y = 16'h200;
			16'h6cf6: y = 16'h200;
			16'h6cf7: y = 16'h200;
			16'h6cf8: y = 16'h200;
			16'h6cf9: y = 16'h200;
			16'h6cfa: y = 16'h200;
			16'h6cfb: y = 16'h200;
			16'h6cfc: y = 16'h200;
			16'h6cfd: y = 16'h200;
			16'h6cfe: y = 16'h200;
			16'h6cff: y = 16'h200;
			16'h6d00: y = 16'h200;
			16'h6d01: y = 16'h200;
			16'h6d02: y = 16'h200;
			16'h6d03: y = 16'h200;
			16'h6d04: y = 16'h200;
			16'h6d05: y = 16'h200;
			16'h6d06: y = 16'h200;
			16'h6d07: y = 16'h200;
			16'h6d08: y = 16'h200;
			16'h6d09: y = 16'h200;
			16'h6d0a: y = 16'h200;
			16'h6d0b: y = 16'h200;
			16'h6d0c: y = 16'h200;
			16'h6d0d: y = 16'h200;
			16'h6d0e: y = 16'h200;
			16'h6d0f: y = 16'h200;
			16'h6d10: y = 16'h200;
			16'h6d11: y = 16'h200;
			16'h6d12: y = 16'h200;
			16'h6d13: y = 16'h200;
			16'h6d14: y = 16'h200;
			16'h6d15: y = 16'h200;
			16'h6d16: y = 16'h200;
			16'h6d17: y = 16'h200;
			16'h6d18: y = 16'h200;
			16'h6d19: y = 16'h200;
			16'h6d1a: y = 16'h200;
			16'h6d1b: y = 16'h200;
			16'h6d1c: y = 16'h200;
			16'h6d1d: y = 16'h200;
			16'h6d1e: y = 16'h200;
			16'h6d1f: y = 16'h200;
			16'h6d20: y = 16'h200;
			16'h6d21: y = 16'h200;
			16'h6d22: y = 16'h200;
			16'h6d23: y = 16'h200;
			16'h6d24: y = 16'h200;
			16'h6d25: y = 16'h200;
			16'h6d26: y = 16'h200;
			16'h6d27: y = 16'h200;
			16'h6d28: y = 16'h200;
			16'h6d29: y = 16'h200;
			16'h6d2a: y = 16'h200;
			16'h6d2b: y = 16'h200;
			16'h6d2c: y = 16'h200;
			16'h6d2d: y = 16'h200;
			16'h6d2e: y = 16'h200;
			16'h6d2f: y = 16'h200;
			16'h6d30: y = 16'h200;
			16'h6d31: y = 16'h200;
			16'h6d32: y = 16'h200;
			16'h6d33: y = 16'h200;
			16'h6d34: y = 16'h200;
			16'h6d35: y = 16'h200;
			16'h6d36: y = 16'h200;
			16'h6d37: y = 16'h200;
			16'h6d38: y = 16'h200;
			16'h6d39: y = 16'h200;
			16'h6d3a: y = 16'h200;
			16'h6d3b: y = 16'h200;
			16'h6d3c: y = 16'h200;
			16'h6d3d: y = 16'h200;
			16'h6d3e: y = 16'h200;
			16'h6d3f: y = 16'h200;
			16'h6d40: y = 16'h200;
			16'h6d41: y = 16'h200;
			16'h6d42: y = 16'h200;
			16'h6d43: y = 16'h200;
			16'h6d44: y = 16'h200;
			16'h6d45: y = 16'h200;
			16'h6d46: y = 16'h200;
			16'h6d47: y = 16'h200;
			16'h6d48: y = 16'h200;
			16'h6d49: y = 16'h200;
			16'h6d4a: y = 16'h200;
			16'h6d4b: y = 16'h200;
			16'h6d4c: y = 16'h200;
			16'h6d4d: y = 16'h200;
			16'h6d4e: y = 16'h200;
			16'h6d4f: y = 16'h200;
			16'h6d50: y = 16'h200;
			16'h6d51: y = 16'h200;
			16'h6d52: y = 16'h200;
			16'h6d53: y = 16'h200;
			16'h6d54: y = 16'h200;
			16'h6d55: y = 16'h200;
			16'h6d56: y = 16'h200;
			16'h6d57: y = 16'h200;
			16'h6d58: y = 16'h200;
			16'h6d59: y = 16'h200;
			16'h6d5a: y = 16'h200;
			16'h6d5b: y = 16'h200;
			16'h6d5c: y = 16'h200;
			16'h6d5d: y = 16'h200;
			16'h6d5e: y = 16'h200;
			16'h6d5f: y = 16'h200;
			16'h6d60: y = 16'h200;
			16'h6d61: y = 16'h200;
			16'h6d62: y = 16'h200;
			16'h6d63: y = 16'h200;
			16'h6d64: y = 16'h200;
			16'h6d65: y = 16'h200;
			16'h6d66: y = 16'h200;
			16'h6d67: y = 16'h200;
			16'h6d68: y = 16'h200;
			16'h6d69: y = 16'h200;
			16'h6d6a: y = 16'h200;
			16'h6d6b: y = 16'h200;
			16'h6d6c: y = 16'h200;
			16'h6d6d: y = 16'h200;
			16'h6d6e: y = 16'h200;
			16'h6d6f: y = 16'h200;
			16'h6d70: y = 16'h200;
			16'h6d71: y = 16'h200;
			16'h6d72: y = 16'h200;
			16'h6d73: y = 16'h200;
			16'h6d74: y = 16'h200;
			16'h6d75: y = 16'h200;
			16'h6d76: y = 16'h200;
			16'h6d77: y = 16'h200;
			16'h6d78: y = 16'h200;
			16'h6d79: y = 16'h200;
			16'h6d7a: y = 16'h200;
			16'h6d7b: y = 16'h200;
			16'h6d7c: y = 16'h200;
			16'h6d7d: y = 16'h200;
			16'h6d7e: y = 16'h200;
			16'h6d7f: y = 16'h200;
			16'h6d80: y = 16'h200;
			16'h6d81: y = 16'h200;
			16'h6d82: y = 16'h200;
			16'h6d83: y = 16'h200;
			16'h6d84: y = 16'h200;
			16'h6d85: y = 16'h200;
			16'h6d86: y = 16'h200;
			16'h6d87: y = 16'h200;
			16'h6d88: y = 16'h200;
			16'h6d89: y = 16'h200;
			16'h6d8a: y = 16'h200;
			16'h6d8b: y = 16'h200;
			16'h6d8c: y = 16'h200;
			16'h6d8d: y = 16'h200;
			16'h6d8e: y = 16'h200;
			16'h6d8f: y = 16'h200;
			16'h6d90: y = 16'h200;
			16'h6d91: y = 16'h200;
			16'h6d92: y = 16'h200;
			16'h6d93: y = 16'h200;
			16'h6d94: y = 16'h200;
			16'h6d95: y = 16'h200;
			16'h6d96: y = 16'h200;
			16'h6d97: y = 16'h200;
			16'h6d98: y = 16'h200;
			16'h6d99: y = 16'h200;
			16'h6d9a: y = 16'h200;
			16'h6d9b: y = 16'h200;
			16'h6d9c: y = 16'h200;
			16'h6d9d: y = 16'h200;
			16'h6d9e: y = 16'h200;
			16'h6d9f: y = 16'h200;
			16'h6da0: y = 16'h200;
			16'h6da1: y = 16'h200;
			16'h6da2: y = 16'h200;
			16'h6da3: y = 16'h200;
			16'h6da4: y = 16'h200;
			16'h6da5: y = 16'h200;
			16'h6da6: y = 16'h200;
			16'h6da7: y = 16'h200;
			16'h6da8: y = 16'h200;
			16'h6da9: y = 16'h200;
			16'h6daa: y = 16'h200;
			16'h6dab: y = 16'h200;
			16'h6dac: y = 16'h200;
			16'h6dad: y = 16'h200;
			16'h6dae: y = 16'h200;
			16'h6daf: y = 16'h200;
			16'h6db0: y = 16'h200;
			16'h6db1: y = 16'h200;
			16'h6db2: y = 16'h200;
			16'h6db3: y = 16'h200;
			16'h6db4: y = 16'h200;
			16'h6db5: y = 16'h200;
			16'h6db6: y = 16'h200;
			16'h6db7: y = 16'h200;
			16'h6db8: y = 16'h200;
			16'h6db9: y = 16'h200;
			16'h6dba: y = 16'h200;
			16'h6dbb: y = 16'h200;
			16'h6dbc: y = 16'h200;
			16'h6dbd: y = 16'h200;
			16'h6dbe: y = 16'h200;
			16'h6dbf: y = 16'h200;
			16'h6dc0: y = 16'h200;
			16'h6dc1: y = 16'h200;
			16'h6dc2: y = 16'h200;
			16'h6dc3: y = 16'h200;
			16'h6dc4: y = 16'h200;
			16'h6dc5: y = 16'h200;
			16'h6dc6: y = 16'h200;
			16'h6dc7: y = 16'h200;
			16'h6dc8: y = 16'h200;
			16'h6dc9: y = 16'h200;
			16'h6dca: y = 16'h200;
			16'h6dcb: y = 16'h200;
			16'h6dcc: y = 16'h200;
			16'h6dcd: y = 16'h200;
			16'h6dce: y = 16'h200;
			16'h6dcf: y = 16'h200;
			16'h6dd0: y = 16'h200;
			16'h6dd1: y = 16'h200;
			16'h6dd2: y = 16'h200;
			16'h6dd3: y = 16'h200;
			16'h6dd4: y = 16'h200;
			16'h6dd5: y = 16'h200;
			16'h6dd6: y = 16'h200;
			16'h6dd7: y = 16'h200;
			16'h6dd8: y = 16'h200;
			16'h6dd9: y = 16'h200;
			16'h6dda: y = 16'h200;
			16'h6ddb: y = 16'h200;
			16'h6ddc: y = 16'h200;
			16'h6ddd: y = 16'h200;
			16'h6dde: y = 16'h200;
			16'h6ddf: y = 16'h200;
			16'h6de0: y = 16'h200;
			16'h6de1: y = 16'h200;
			16'h6de2: y = 16'h200;
			16'h6de3: y = 16'h200;
			16'h6de4: y = 16'h200;
			16'h6de5: y = 16'h200;
			16'h6de6: y = 16'h200;
			16'h6de7: y = 16'h200;
			16'h6de8: y = 16'h200;
			16'h6de9: y = 16'h200;
			16'h6dea: y = 16'h200;
			16'h6deb: y = 16'h200;
			16'h6dec: y = 16'h200;
			16'h6ded: y = 16'h200;
			16'h6dee: y = 16'h200;
			16'h6def: y = 16'h200;
			16'h6df0: y = 16'h200;
			16'h6df1: y = 16'h200;
			16'h6df2: y = 16'h200;
			16'h6df3: y = 16'h200;
			16'h6df4: y = 16'h200;
			16'h6df5: y = 16'h200;
			16'h6df6: y = 16'h200;
			16'h6df7: y = 16'h200;
			16'h6df8: y = 16'h200;
			16'h6df9: y = 16'h200;
			16'h6dfa: y = 16'h200;
			16'h6dfb: y = 16'h200;
			16'h6dfc: y = 16'h200;
			16'h6dfd: y = 16'h200;
			16'h6dfe: y = 16'h200;
			16'h6dff: y = 16'h200;
			16'h6e00: y = 16'h200;
			16'h6e01: y = 16'h200;
			16'h6e02: y = 16'h200;
			16'h6e03: y = 16'h200;
			16'h6e04: y = 16'h200;
			16'h6e05: y = 16'h200;
			16'h6e06: y = 16'h200;
			16'h6e07: y = 16'h200;
			16'h6e08: y = 16'h200;
			16'h6e09: y = 16'h200;
			16'h6e0a: y = 16'h200;
			16'h6e0b: y = 16'h200;
			16'h6e0c: y = 16'h200;
			16'h6e0d: y = 16'h200;
			16'h6e0e: y = 16'h200;
			16'h6e0f: y = 16'h200;
			16'h6e10: y = 16'h200;
			16'h6e11: y = 16'h200;
			16'h6e12: y = 16'h200;
			16'h6e13: y = 16'h200;
			16'h6e14: y = 16'h200;
			16'h6e15: y = 16'h200;
			16'h6e16: y = 16'h200;
			16'h6e17: y = 16'h200;
			16'h6e18: y = 16'h200;
			16'h6e19: y = 16'h200;
			16'h6e1a: y = 16'h200;
			16'h6e1b: y = 16'h200;
			16'h6e1c: y = 16'h200;
			16'h6e1d: y = 16'h200;
			16'h6e1e: y = 16'h200;
			16'h6e1f: y = 16'h200;
			16'h6e20: y = 16'h200;
			16'h6e21: y = 16'h200;
			16'h6e22: y = 16'h200;
			16'h6e23: y = 16'h200;
			16'h6e24: y = 16'h200;
			16'h6e25: y = 16'h200;
			16'h6e26: y = 16'h200;
			16'h6e27: y = 16'h200;
			16'h6e28: y = 16'h200;
			16'h6e29: y = 16'h200;
			16'h6e2a: y = 16'h200;
			16'h6e2b: y = 16'h200;
			16'h6e2c: y = 16'h200;
			16'h6e2d: y = 16'h200;
			16'h6e2e: y = 16'h200;
			16'h6e2f: y = 16'h200;
			16'h6e30: y = 16'h200;
			16'h6e31: y = 16'h200;
			16'h6e32: y = 16'h200;
			16'h6e33: y = 16'h200;
			16'h6e34: y = 16'h200;
			16'h6e35: y = 16'h200;
			16'h6e36: y = 16'h200;
			16'h6e37: y = 16'h200;
			16'h6e38: y = 16'h200;
			16'h6e39: y = 16'h200;
			16'h6e3a: y = 16'h200;
			16'h6e3b: y = 16'h200;
			16'h6e3c: y = 16'h200;
			16'h6e3d: y = 16'h200;
			16'h6e3e: y = 16'h200;
			16'h6e3f: y = 16'h200;
			16'h6e40: y = 16'h200;
			16'h6e41: y = 16'h200;
			16'h6e42: y = 16'h200;
			16'h6e43: y = 16'h200;
			16'h6e44: y = 16'h200;
			16'h6e45: y = 16'h200;
			16'h6e46: y = 16'h200;
			16'h6e47: y = 16'h200;
			16'h6e48: y = 16'h200;
			16'h6e49: y = 16'h200;
			16'h6e4a: y = 16'h200;
			16'h6e4b: y = 16'h200;
			16'h6e4c: y = 16'h200;
			16'h6e4d: y = 16'h200;
			16'h6e4e: y = 16'h200;
			16'h6e4f: y = 16'h200;
			16'h6e50: y = 16'h200;
			16'h6e51: y = 16'h200;
			16'h6e52: y = 16'h200;
			16'h6e53: y = 16'h200;
			16'h6e54: y = 16'h200;
			16'h6e55: y = 16'h200;
			16'h6e56: y = 16'h200;
			16'h6e57: y = 16'h200;
			16'h6e58: y = 16'h200;
			16'h6e59: y = 16'h200;
			16'h6e5a: y = 16'h200;
			16'h6e5b: y = 16'h200;
			16'h6e5c: y = 16'h200;
			16'h6e5d: y = 16'h200;
			16'h6e5e: y = 16'h200;
			16'h6e5f: y = 16'h200;
			16'h6e60: y = 16'h200;
			16'h6e61: y = 16'h200;
			16'h6e62: y = 16'h200;
			16'h6e63: y = 16'h200;
			16'h6e64: y = 16'h200;
			16'h6e65: y = 16'h200;
			16'h6e66: y = 16'h200;
			16'h6e67: y = 16'h200;
			16'h6e68: y = 16'h200;
			16'h6e69: y = 16'h200;
			16'h6e6a: y = 16'h200;
			16'h6e6b: y = 16'h200;
			16'h6e6c: y = 16'h200;
			16'h6e6d: y = 16'h200;
			16'h6e6e: y = 16'h200;
			16'h6e6f: y = 16'h200;
			16'h6e70: y = 16'h200;
			16'h6e71: y = 16'h200;
			16'h6e72: y = 16'h200;
			16'h6e73: y = 16'h200;
			16'h6e74: y = 16'h200;
			16'h6e75: y = 16'h200;
			16'h6e76: y = 16'h200;
			16'h6e77: y = 16'h200;
			16'h6e78: y = 16'h200;
			16'h6e79: y = 16'h200;
			16'h6e7a: y = 16'h200;
			16'h6e7b: y = 16'h200;
			16'h6e7c: y = 16'h200;
			16'h6e7d: y = 16'h200;
			16'h6e7e: y = 16'h200;
			16'h6e7f: y = 16'h200;
			16'h6e80: y = 16'h200;
			16'h6e81: y = 16'h200;
			16'h6e82: y = 16'h200;
			16'h6e83: y = 16'h200;
			16'h6e84: y = 16'h200;
			16'h6e85: y = 16'h200;
			16'h6e86: y = 16'h200;
			16'h6e87: y = 16'h200;
			16'h6e88: y = 16'h200;
			16'h6e89: y = 16'h200;
			16'h6e8a: y = 16'h200;
			16'h6e8b: y = 16'h200;
			16'h6e8c: y = 16'h200;
			16'h6e8d: y = 16'h200;
			16'h6e8e: y = 16'h200;
			16'h6e8f: y = 16'h200;
			16'h6e90: y = 16'h200;
			16'h6e91: y = 16'h200;
			16'h6e92: y = 16'h200;
			16'h6e93: y = 16'h200;
			16'h6e94: y = 16'h200;
			16'h6e95: y = 16'h200;
			16'h6e96: y = 16'h200;
			16'h6e97: y = 16'h200;
			16'h6e98: y = 16'h200;
			16'h6e99: y = 16'h200;
			16'h6e9a: y = 16'h200;
			16'h6e9b: y = 16'h200;
			16'h6e9c: y = 16'h200;
			16'h6e9d: y = 16'h200;
			16'h6e9e: y = 16'h200;
			16'h6e9f: y = 16'h200;
			16'h6ea0: y = 16'h200;
			16'h6ea1: y = 16'h200;
			16'h6ea2: y = 16'h200;
			16'h6ea3: y = 16'h200;
			16'h6ea4: y = 16'h200;
			16'h6ea5: y = 16'h200;
			16'h6ea6: y = 16'h200;
			16'h6ea7: y = 16'h200;
			16'h6ea8: y = 16'h200;
			16'h6ea9: y = 16'h200;
			16'h6eaa: y = 16'h200;
			16'h6eab: y = 16'h200;
			16'h6eac: y = 16'h200;
			16'h6ead: y = 16'h200;
			16'h6eae: y = 16'h200;
			16'h6eaf: y = 16'h200;
			16'h6eb0: y = 16'h200;
			16'h6eb1: y = 16'h200;
			16'h6eb2: y = 16'h200;
			16'h6eb3: y = 16'h200;
			16'h6eb4: y = 16'h200;
			16'h6eb5: y = 16'h200;
			16'h6eb6: y = 16'h200;
			16'h6eb7: y = 16'h200;
			16'h6eb8: y = 16'h200;
			16'h6eb9: y = 16'h200;
			16'h6eba: y = 16'h200;
			16'h6ebb: y = 16'h200;
			16'h6ebc: y = 16'h200;
			16'h6ebd: y = 16'h200;
			16'h6ebe: y = 16'h200;
			16'h6ebf: y = 16'h200;
			16'h6ec0: y = 16'h200;
			16'h6ec1: y = 16'h200;
			16'h6ec2: y = 16'h200;
			16'h6ec3: y = 16'h200;
			16'h6ec4: y = 16'h200;
			16'h6ec5: y = 16'h200;
			16'h6ec6: y = 16'h200;
			16'h6ec7: y = 16'h200;
			16'h6ec8: y = 16'h200;
			16'h6ec9: y = 16'h200;
			16'h6eca: y = 16'h200;
			16'h6ecb: y = 16'h200;
			16'h6ecc: y = 16'h200;
			16'h6ecd: y = 16'h200;
			16'h6ece: y = 16'h200;
			16'h6ecf: y = 16'h200;
			16'h6ed0: y = 16'h200;
			16'h6ed1: y = 16'h200;
			16'h6ed2: y = 16'h200;
			16'h6ed3: y = 16'h200;
			16'h6ed4: y = 16'h200;
			16'h6ed5: y = 16'h200;
			16'h6ed6: y = 16'h200;
			16'h6ed7: y = 16'h200;
			16'h6ed8: y = 16'h200;
			16'h6ed9: y = 16'h200;
			16'h6eda: y = 16'h200;
			16'h6edb: y = 16'h200;
			16'h6edc: y = 16'h200;
			16'h6edd: y = 16'h200;
			16'h6ede: y = 16'h200;
			16'h6edf: y = 16'h200;
			16'h6ee0: y = 16'h200;
			16'h6ee1: y = 16'h200;
			16'h6ee2: y = 16'h200;
			16'h6ee3: y = 16'h200;
			16'h6ee4: y = 16'h200;
			16'h6ee5: y = 16'h200;
			16'h6ee6: y = 16'h200;
			16'h6ee7: y = 16'h200;
			16'h6ee8: y = 16'h200;
			16'h6ee9: y = 16'h200;
			16'h6eea: y = 16'h200;
			16'h6eeb: y = 16'h200;
			16'h6eec: y = 16'h200;
			16'h6eed: y = 16'h200;
			16'h6eee: y = 16'h200;
			16'h6eef: y = 16'h200;
			16'h6ef0: y = 16'h200;
			16'h6ef1: y = 16'h200;
			16'h6ef2: y = 16'h200;
			16'h6ef3: y = 16'h200;
			16'h6ef4: y = 16'h200;
			16'h6ef5: y = 16'h200;
			16'h6ef6: y = 16'h200;
			16'h6ef7: y = 16'h200;
			16'h6ef8: y = 16'h200;
			16'h6ef9: y = 16'h200;
			16'h6efa: y = 16'h200;
			16'h6efb: y = 16'h200;
			16'h6efc: y = 16'h200;
			16'h6efd: y = 16'h200;
			16'h6efe: y = 16'h200;
			16'h6eff: y = 16'h200;
			16'h6f00: y = 16'h200;
			16'h6f01: y = 16'h200;
			16'h6f02: y = 16'h200;
			16'h6f03: y = 16'h200;
			16'h6f04: y = 16'h200;
			16'h6f05: y = 16'h200;
			16'h6f06: y = 16'h200;
			16'h6f07: y = 16'h200;
			16'h6f08: y = 16'h200;
			16'h6f09: y = 16'h200;
			16'h6f0a: y = 16'h200;
			16'h6f0b: y = 16'h200;
			16'h6f0c: y = 16'h200;
			16'h6f0d: y = 16'h200;
			16'h6f0e: y = 16'h200;
			16'h6f0f: y = 16'h200;
			16'h6f10: y = 16'h200;
			16'h6f11: y = 16'h200;
			16'h6f12: y = 16'h200;
			16'h6f13: y = 16'h200;
			16'h6f14: y = 16'h200;
			16'h6f15: y = 16'h200;
			16'h6f16: y = 16'h200;
			16'h6f17: y = 16'h200;
			16'h6f18: y = 16'h200;
			16'h6f19: y = 16'h200;
			16'h6f1a: y = 16'h200;
			16'h6f1b: y = 16'h200;
			16'h6f1c: y = 16'h200;
			16'h6f1d: y = 16'h200;
			16'h6f1e: y = 16'h200;
			16'h6f1f: y = 16'h200;
			16'h6f20: y = 16'h200;
			16'h6f21: y = 16'h200;
			16'h6f22: y = 16'h200;
			16'h6f23: y = 16'h200;
			16'h6f24: y = 16'h200;
			16'h6f25: y = 16'h200;
			16'h6f26: y = 16'h200;
			16'h6f27: y = 16'h200;
			16'h6f28: y = 16'h200;
			16'h6f29: y = 16'h200;
			16'h6f2a: y = 16'h200;
			16'h6f2b: y = 16'h200;
			16'h6f2c: y = 16'h200;
			16'h6f2d: y = 16'h200;
			16'h6f2e: y = 16'h200;
			16'h6f2f: y = 16'h200;
			16'h6f30: y = 16'h200;
			16'h6f31: y = 16'h200;
			16'h6f32: y = 16'h200;
			16'h6f33: y = 16'h200;
			16'h6f34: y = 16'h200;
			16'h6f35: y = 16'h200;
			16'h6f36: y = 16'h200;
			16'h6f37: y = 16'h200;
			16'h6f38: y = 16'h200;
			16'h6f39: y = 16'h200;
			16'h6f3a: y = 16'h200;
			16'h6f3b: y = 16'h200;
			16'h6f3c: y = 16'h200;
			16'h6f3d: y = 16'h200;
			16'h6f3e: y = 16'h200;
			16'h6f3f: y = 16'h200;
			16'h6f40: y = 16'h200;
			16'h6f41: y = 16'h200;
			16'h6f42: y = 16'h200;
			16'h6f43: y = 16'h200;
			16'h6f44: y = 16'h200;
			16'h6f45: y = 16'h200;
			16'h6f46: y = 16'h200;
			16'h6f47: y = 16'h200;
			16'h6f48: y = 16'h200;
			16'h6f49: y = 16'h200;
			16'h6f4a: y = 16'h200;
			16'h6f4b: y = 16'h200;
			16'h6f4c: y = 16'h200;
			16'h6f4d: y = 16'h200;
			16'h6f4e: y = 16'h200;
			16'h6f4f: y = 16'h200;
			16'h6f50: y = 16'h200;
			16'h6f51: y = 16'h200;
			16'h6f52: y = 16'h200;
			16'h6f53: y = 16'h200;
			16'h6f54: y = 16'h200;
			16'h6f55: y = 16'h200;
			16'h6f56: y = 16'h200;
			16'h6f57: y = 16'h200;
			16'h6f58: y = 16'h200;
			16'h6f59: y = 16'h200;
			16'h6f5a: y = 16'h200;
			16'h6f5b: y = 16'h200;
			16'h6f5c: y = 16'h200;
			16'h6f5d: y = 16'h200;
			16'h6f5e: y = 16'h200;
			16'h6f5f: y = 16'h200;
			16'h6f60: y = 16'h200;
			16'h6f61: y = 16'h200;
			16'h6f62: y = 16'h200;
			16'h6f63: y = 16'h200;
			16'h6f64: y = 16'h200;
			16'h6f65: y = 16'h200;
			16'h6f66: y = 16'h200;
			16'h6f67: y = 16'h200;
			16'h6f68: y = 16'h200;
			16'h6f69: y = 16'h200;
			16'h6f6a: y = 16'h200;
			16'h6f6b: y = 16'h200;
			16'h6f6c: y = 16'h200;
			16'h6f6d: y = 16'h200;
			16'h6f6e: y = 16'h200;
			16'h6f6f: y = 16'h200;
			16'h6f70: y = 16'h200;
			16'h6f71: y = 16'h200;
			16'h6f72: y = 16'h200;
			16'h6f73: y = 16'h200;
			16'h6f74: y = 16'h200;
			16'h6f75: y = 16'h200;
			16'h6f76: y = 16'h200;
			16'h6f77: y = 16'h200;
			16'h6f78: y = 16'h200;
			16'h6f79: y = 16'h200;
			16'h6f7a: y = 16'h200;
			16'h6f7b: y = 16'h200;
			16'h6f7c: y = 16'h200;
			16'h6f7d: y = 16'h200;
			16'h6f7e: y = 16'h200;
			16'h6f7f: y = 16'h200;
			16'h6f80: y = 16'h200;
			16'h6f81: y = 16'h200;
			16'h6f82: y = 16'h200;
			16'h6f83: y = 16'h200;
			16'h6f84: y = 16'h200;
			16'h6f85: y = 16'h200;
			16'h6f86: y = 16'h200;
			16'h6f87: y = 16'h200;
			16'h6f88: y = 16'h200;
			16'h6f89: y = 16'h200;
			16'h6f8a: y = 16'h200;
			16'h6f8b: y = 16'h200;
			16'h6f8c: y = 16'h200;
			16'h6f8d: y = 16'h200;
			16'h6f8e: y = 16'h200;
			16'h6f8f: y = 16'h200;
			16'h6f90: y = 16'h200;
			16'h6f91: y = 16'h200;
			16'h6f92: y = 16'h200;
			16'h6f93: y = 16'h200;
			16'h6f94: y = 16'h200;
			16'h6f95: y = 16'h200;
			16'h6f96: y = 16'h200;
			16'h6f97: y = 16'h200;
			16'h6f98: y = 16'h200;
			16'h6f99: y = 16'h200;
			16'h6f9a: y = 16'h200;
			16'h6f9b: y = 16'h200;
			16'h6f9c: y = 16'h200;
			16'h6f9d: y = 16'h200;
			16'h6f9e: y = 16'h200;
			16'h6f9f: y = 16'h200;
			16'h6fa0: y = 16'h200;
			16'h6fa1: y = 16'h200;
			16'h6fa2: y = 16'h200;
			16'h6fa3: y = 16'h200;
			16'h6fa4: y = 16'h200;
			16'h6fa5: y = 16'h200;
			16'h6fa6: y = 16'h200;
			16'h6fa7: y = 16'h200;
			16'h6fa8: y = 16'h200;
			16'h6fa9: y = 16'h200;
			16'h6faa: y = 16'h200;
			16'h6fab: y = 16'h200;
			16'h6fac: y = 16'h200;
			16'h6fad: y = 16'h200;
			16'h6fae: y = 16'h200;
			16'h6faf: y = 16'h200;
			16'h6fb0: y = 16'h200;
			16'h6fb1: y = 16'h200;
			16'h6fb2: y = 16'h200;
			16'h6fb3: y = 16'h200;
			16'h6fb4: y = 16'h200;
			16'h6fb5: y = 16'h200;
			16'h6fb6: y = 16'h200;
			16'h6fb7: y = 16'h200;
			16'h6fb8: y = 16'h200;
			16'h6fb9: y = 16'h200;
			16'h6fba: y = 16'h200;
			16'h6fbb: y = 16'h200;
			16'h6fbc: y = 16'h200;
			16'h6fbd: y = 16'h200;
			16'h6fbe: y = 16'h200;
			16'h6fbf: y = 16'h200;
			16'h6fc0: y = 16'h200;
			16'h6fc1: y = 16'h200;
			16'h6fc2: y = 16'h200;
			16'h6fc3: y = 16'h200;
			16'h6fc4: y = 16'h200;
			16'h6fc5: y = 16'h200;
			16'h6fc6: y = 16'h200;
			16'h6fc7: y = 16'h200;
			16'h6fc8: y = 16'h200;
			16'h6fc9: y = 16'h200;
			16'h6fca: y = 16'h200;
			16'h6fcb: y = 16'h200;
			16'h6fcc: y = 16'h200;
			16'h6fcd: y = 16'h200;
			16'h6fce: y = 16'h200;
			16'h6fcf: y = 16'h200;
			16'h6fd0: y = 16'h200;
			16'h6fd1: y = 16'h200;
			16'h6fd2: y = 16'h200;
			16'h6fd3: y = 16'h200;
			16'h6fd4: y = 16'h200;
			16'h6fd5: y = 16'h200;
			16'h6fd6: y = 16'h200;
			16'h6fd7: y = 16'h200;
			16'h6fd8: y = 16'h200;
			16'h6fd9: y = 16'h200;
			16'h6fda: y = 16'h200;
			16'h6fdb: y = 16'h200;
			16'h6fdc: y = 16'h200;
			16'h6fdd: y = 16'h200;
			16'h6fde: y = 16'h200;
			16'h6fdf: y = 16'h200;
			16'h6fe0: y = 16'h200;
			16'h6fe1: y = 16'h200;
			16'h6fe2: y = 16'h200;
			16'h6fe3: y = 16'h200;
			16'h6fe4: y = 16'h200;
			16'h6fe5: y = 16'h200;
			16'h6fe6: y = 16'h200;
			16'h6fe7: y = 16'h200;
			16'h6fe8: y = 16'h200;
			16'h6fe9: y = 16'h200;
			16'h6fea: y = 16'h200;
			16'h6feb: y = 16'h200;
			16'h6fec: y = 16'h200;
			16'h6fed: y = 16'h200;
			16'h6fee: y = 16'h200;
			16'h6fef: y = 16'h200;
			16'h6ff0: y = 16'h200;
			16'h6ff1: y = 16'h200;
			16'h6ff2: y = 16'h200;
			16'h6ff3: y = 16'h200;
			16'h6ff4: y = 16'h200;
			16'h6ff5: y = 16'h200;
			16'h6ff6: y = 16'h200;
			16'h6ff7: y = 16'h200;
			16'h6ff8: y = 16'h200;
			16'h6ff9: y = 16'h200;
			16'h6ffa: y = 16'h200;
			16'h6ffb: y = 16'h200;
			16'h6ffc: y = 16'h200;
			16'h6ffd: y = 16'h200;
			16'h6ffe: y = 16'h200;
			16'h6fff: y = 16'h200;
			16'h7000: y = 16'h200;
			16'h7001: y = 16'h200;
			16'h7002: y = 16'h200;
			16'h7003: y = 16'h200;
			16'h7004: y = 16'h200;
			16'h7005: y = 16'h200;
			16'h7006: y = 16'h200;
			16'h7007: y = 16'h200;
			16'h7008: y = 16'h200;
			16'h7009: y = 16'h200;
			16'h700a: y = 16'h200;
			16'h700b: y = 16'h200;
			16'h700c: y = 16'h200;
			16'h700d: y = 16'h200;
			16'h700e: y = 16'h200;
			16'h700f: y = 16'h200;
			16'h7010: y = 16'h200;
			16'h7011: y = 16'h200;
			16'h7012: y = 16'h200;
			16'h7013: y = 16'h200;
			16'h7014: y = 16'h200;
			16'h7015: y = 16'h200;
			16'h7016: y = 16'h200;
			16'h7017: y = 16'h200;
			16'h7018: y = 16'h200;
			16'h7019: y = 16'h200;
			16'h701a: y = 16'h200;
			16'h701b: y = 16'h200;
			16'h701c: y = 16'h200;
			16'h701d: y = 16'h200;
			16'h701e: y = 16'h200;
			16'h701f: y = 16'h200;
			16'h7020: y = 16'h200;
			16'h7021: y = 16'h200;
			16'h7022: y = 16'h200;
			16'h7023: y = 16'h200;
			16'h7024: y = 16'h200;
			16'h7025: y = 16'h200;
			16'h7026: y = 16'h200;
			16'h7027: y = 16'h200;
			16'h7028: y = 16'h200;
			16'h7029: y = 16'h200;
			16'h702a: y = 16'h200;
			16'h702b: y = 16'h200;
			16'h702c: y = 16'h200;
			16'h702d: y = 16'h200;
			16'h702e: y = 16'h200;
			16'h702f: y = 16'h200;
			16'h7030: y = 16'h200;
			16'h7031: y = 16'h200;
			16'h7032: y = 16'h200;
			16'h7033: y = 16'h200;
			16'h7034: y = 16'h200;
			16'h7035: y = 16'h200;
			16'h7036: y = 16'h200;
			16'h7037: y = 16'h200;
			16'h7038: y = 16'h200;
			16'h7039: y = 16'h200;
			16'h703a: y = 16'h200;
			16'h703b: y = 16'h200;
			16'h703c: y = 16'h200;
			16'h703d: y = 16'h200;
			16'h703e: y = 16'h200;
			16'h703f: y = 16'h200;
			16'h7040: y = 16'h200;
			16'h7041: y = 16'h200;
			16'h7042: y = 16'h200;
			16'h7043: y = 16'h200;
			16'h7044: y = 16'h200;
			16'h7045: y = 16'h200;
			16'h7046: y = 16'h200;
			16'h7047: y = 16'h200;
			16'h7048: y = 16'h200;
			16'h7049: y = 16'h200;
			16'h704a: y = 16'h200;
			16'h704b: y = 16'h200;
			16'h704c: y = 16'h200;
			16'h704d: y = 16'h200;
			16'h704e: y = 16'h200;
			16'h704f: y = 16'h200;
			16'h7050: y = 16'h200;
			16'h7051: y = 16'h200;
			16'h7052: y = 16'h200;
			16'h7053: y = 16'h200;
			16'h7054: y = 16'h200;
			16'h7055: y = 16'h200;
			16'h7056: y = 16'h200;
			16'h7057: y = 16'h200;
			16'h7058: y = 16'h200;
			16'h7059: y = 16'h200;
			16'h705a: y = 16'h200;
			16'h705b: y = 16'h200;
			16'h705c: y = 16'h200;
			16'h705d: y = 16'h200;
			16'h705e: y = 16'h200;
			16'h705f: y = 16'h200;
			16'h7060: y = 16'h200;
			16'h7061: y = 16'h200;
			16'h7062: y = 16'h200;
			16'h7063: y = 16'h200;
			16'h7064: y = 16'h200;
			16'h7065: y = 16'h200;
			16'h7066: y = 16'h200;
			16'h7067: y = 16'h200;
			16'h7068: y = 16'h200;
			16'h7069: y = 16'h200;
			16'h706a: y = 16'h200;
			16'h706b: y = 16'h200;
			16'h706c: y = 16'h200;
			16'h706d: y = 16'h200;
			16'h706e: y = 16'h200;
			16'h706f: y = 16'h200;
			16'h7070: y = 16'h200;
			16'h7071: y = 16'h200;
			16'h7072: y = 16'h200;
			16'h7073: y = 16'h200;
			16'h7074: y = 16'h200;
			16'h7075: y = 16'h200;
			16'h7076: y = 16'h200;
			16'h7077: y = 16'h200;
			16'h7078: y = 16'h200;
			16'h7079: y = 16'h200;
			16'h707a: y = 16'h200;
			16'h707b: y = 16'h200;
			16'h707c: y = 16'h200;
			16'h707d: y = 16'h200;
			16'h707e: y = 16'h200;
			16'h707f: y = 16'h200;
			16'h7080: y = 16'h200;
			16'h7081: y = 16'h200;
			16'h7082: y = 16'h200;
			16'h7083: y = 16'h200;
			16'h7084: y = 16'h200;
			16'h7085: y = 16'h200;
			16'h7086: y = 16'h200;
			16'h7087: y = 16'h200;
			16'h7088: y = 16'h200;
			16'h7089: y = 16'h200;
			16'h708a: y = 16'h200;
			16'h708b: y = 16'h200;
			16'h708c: y = 16'h200;
			16'h708d: y = 16'h200;
			16'h708e: y = 16'h200;
			16'h708f: y = 16'h200;
			16'h7090: y = 16'h200;
			16'h7091: y = 16'h200;
			16'h7092: y = 16'h200;
			16'h7093: y = 16'h200;
			16'h7094: y = 16'h200;
			16'h7095: y = 16'h200;
			16'h7096: y = 16'h200;
			16'h7097: y = 16'h200;
			16'h7098: y = 16'h200;
			16'h7099: y = 16'h200;
			16'h709a: y = 16'h200;
			16'h709b: y = 16'h200;
			16'h709c: y = 16'h200;
			16'h709d: y = 16'h200;
			16'h709e: y = 16'h200;
			16'h709f: y = 16'h200;
			16'h70a0: y = 16'h200;
			16'h70a1: y = 16'h200;
			16'h70a2: y = 16'h200;
			16'h70a3: y = 16'h200;
			16'h70a4: y = 16'h200;
			16'h70a5: y = 16'h200;
			16'h70a6: y = 16'h200;
			16'h70a7: y = 16'h200;
			16'h70a8: y = 16'h200;
			16'h70a9: y = 16'h200;
			16'h70aa: y = 16'h200;
			16'h70ab: y = 16'h200;
			16'h70ac: y = 16'h200;
			16'h70ad: y = 16'h200;
			16'h70ae: y = 16'h200;
			16'h70af: y = 16'h200;
			16'h70b0: y = 16'h200;
			16'h70b1: y = 16'h200;
			16'h70b2: y = 16'h200;
			16'h70b3: y = 16'h200;
			16'h70b4: y = 16'h200;
			16'h70b5: y = 16'h200;
			16'h70b6: y = 16'h200;
			16'h70b7: y = 16'h200;
			16'h70b8: y = 16'h200;
			16'h70b9: y = 16'h200;
			16'h70ba: y = 16'h200;
			16'h70bb: y = 16'h200;
			16'h70bc: y = 16'h200;
			16'h70bd: y = 16'h200;
			16'h70be: y = 16'h200;
			16'h70bf: y = 16'h200;
			16'h70c0: y = 16'h200;
			16'h70c1: y = 16'h200;
			16'h70c2: y = 16'h200;
			16'h70c3: y = 16'h200;
			16'h70c4: y = 16'h200;
			16'h70c5: y = 16'h200;
			16'h70c6: y = 16'h200;
			16'h70c7: y = 16'h200;
			16'h70c8: y = 16'h200;
			16'h70c9: y = 16'h200;
			16'h70ca: y = 16'h200;
			16'h70cb: y = 16'h200;
			16'h70cc: y = 16'h200;
			16'h70cd: y = 16'h200;
			16'h70ce: y = 16'h200;
			16'h70cf: y = 16'h200;
			16'h70d0: y = 16'h200;
			16'h70d1: y = 16'h200;
			16'h70d2: y = 16'h200;
			16'h70d3: y = 16'h200;
			16'h70d4: y = 16'h200;
			16'h70d5: y = 16'h200;
			16'h70d6: y = 16'h200;
			16'h70d7: y = 16'h200;
			16'h70d8: y = 16'h200;
			16'h70d9: y = 16'h200;
			16'h70da: y = 16'h200;
			16'h70db: y = 16'h200;
			16'h70dc: y = 16'h200;
			16'h70dd: y = 16'h200;
			16'h70de: y = 16'h200;
			16'h70df: y = 16'h200;
			16'h70e0: y = 16'h200;
			16'h70e1: y = 16'h200;
			16'h70e2: y = 16'h200;
			16'h70e3: y = 16'h200;
			16'h70e4: y = 16'h200;
			16'h70e5: y = 16'h200;
			16'h70e6: y = 16'h200;
			16'h70e7: y = 16'h200;
			16'h70e8: y = 16'h200;
			16'h70e9: y = 16'h200;
			16'h70ea: y = 16'h200;
			16'h70eb: y = 16'h200;
			16'h70ec: y = 16'h200;
			16'h70ed: y = 16'h200;
			16'h70ee: y = 16'h200;
			16'h70ef: y = 16'h200;
			16'h70f0: y = 16'h200;
			16'h70f1: y = 16'h200;
			16'h70f2: y = 16'h200;
			16'h70f3: y = 16'h200;
			16'h70f4: y = 16'h200;
			16'h70f5: y = 16'h200;
			16'h70f6: y = 16'h200;
			16'h70f7: y = 16'h200;
			16'h70f8: y = 16'h200;
			16'h70f9: y = 16'h200;
			16'h70fa: y = 16'h200;
			16'h70fb: y = 16'h200;
			16'h70fc: y = 16'h200;
			16'h70fd: y = 16'h200;
			16'h70fe: y = 16'h200;
			16'h70ff: y = 16'h200;
			16'h7100: y = 16'h200;
			16'h7101: y = 16'h200;
			16'h7102: y = 16'h200;
			16'h7103: y = 16'h200;
			16'h7104: y = 16'h200;
			16'h7105: y = 16'h200;
			16'h7106: y = 16'h200;
			16'h7107: y = 16'h200;
			16'h7108: y = 16'h200;
			16'h7109: y = 16'h200;
			16'h710a: y = 16'h200;
			16'h710b: y = 16'h200;
			16'h710c: y = 16'h200;
			16'h710d: y = 16'h200;
			16'h710e: y = 16'h200;
			16'h710f: y = 16'h200;
			16'h7110: y = 16'h200;
			16'h7111: y = 16'h200;
			16'h7112: y = 16'h200;
			16'h7113: y = 16'h200;
			16'h7114: y = 16'h200;
			16'h7115: y = 16'h200;
			16'h7116: y = 16'h200;
			16'h7117: y = 16'h200;
			16'h7118: y = 16'h200;
			16'h7119: y = 16'h200;
			16'h711a: y = 16'h200;
			16'h711b: y = 16'h200;
			16'h711c: y = 16'h200;
			16'h711d: y = 16'h200;
			16'h711e: y = 16'h200;
			16'h711f: y = 16'h200;
			16'h7120: y = 16'h200;
			16'h7121: y = 16'h200;
			16'h7122: y = 16'h200;
			16'h7123: y = 16'h200;
			16'h7124: y = 16'h200;
			16'h7125: y = 16'h200;
			16'h7126: y = 16'h200;
			16'h7127: y = 16'h200;
			16'h7128: y = 16'h200;
			16'h7129: y = 16'h200;
			16'h712a: y = 16'h200;
			16'h712b: y = 16'h200;
			16'h712c: y = 16'h200;
			16'h712d: y = 16'h200;
			16'h712e: y = 16'h200;
			16'h712f: y = 16'h200;
			16'h7130: y = 16'h200;
			16'h7131: y = 16'h200;
			16'h7132: y = 16'h200;
			16'h7133: y = 16'h200;
			16'h7134: y = 16'h200;
			16'h7135: y = 16'h200;
			16'h7136: y = 16'h200;
			16'h7137: y = 16'h200;
			16'h7138: y = 16'h200;
			16'h7139: y = 16'h200;
			16'h713a: y = 16'h200;
			16'h713b: y = 16'h200;
			16'h713c: y = 16'h200;
			16'h713d: y = 16'h200;
			16'h713e: y = 16'h200;
			16'h713f: y = 16'h200;
			16'h7140: y = 16'h200;
			16'h7141: y = 16'h200;
			16'h7142: y = 16'h200;
			16'h7143: y = 16'h200;
			16'h7144: y = 16'h200;
			16'h7145: y = 16'h200;
			16'h7146: y = 16'h200;
			16'h7147: y = 16'h200;
			16'h7148: y = 16'h200;
			16'h7149: y = 16'h200;
			16'h714a: y = 16'h200;
			16'h714b: y = 16'h200;
			16'h714c: y = 16'h200;
			16'h714d: y = 16'h200;
			16'h714e: y = 16'h200;
			16'h714f: y = 16'h200;
			16'h7150: y = 16'h200;
			16'h7151: y = 16'h200;
			16'h7152: y = 16'h200;
			16'h7153: y = 16'h200;
			16'h7154: y = 16'h200;
			16'h7155: y = 16'h200;
			16'h7156: y = 16'h200;
			16'h7157: y = 16'h200;
			16'h7158: y = 16'h200;
			16'h7159: y = 16'h200;
			16'h715a: y = 16'h200;
			16'h715b: y = 16'h200;
			16'h715c: y = 16'h200;
			16'h715d: y = 16'h200;
			16'h715e: y = 16'h200;
			16'h715f: y = 16'h200;
			16'h7160: y = 16'h200;
			16'h7161: y = 16'h200;
			16'h7162: y = 16'h200;
			16'h7163: y = 16'h200;
			16'h7164: y = 16'h200;
			16'h7165: y = 16'h200;
			16'h7166: y = 16'h200;
			16'h7167: y = 16'h200;
			16'h7168: y = 16'h200;
			16'h7169: y = 16'h200;
			16'h716a: y = 16'h200;
			16'h716b: y = 16'h200;
			16'h716c: y = 16'h200;
			16'h716d: y = 16'h200;
			16'h716e: y = 16'h200;
			16'h716f: y = 16'h200;
			16'h7170: y = 16'h200;
			16'h7171: y = 16'h200;
			16'h7172: y = 16'h200;
			16'h7173: y = 16'h200;
			16'h7174: y = 16'h200;
			16'h7175: y = 16'h200;
			16'h7176: y = 16'h200;
			16'h7177: y = 16'h200;
			16'h7178: y = 16'h200;
			16'h7179: y = 16'h200;
			16'h717a: y = 16'h200;
			16'h717b: y = 16'h200;
			16'h717c: y = 16'h200;
			16'h717d: y = 16'h200;
			16'h717e: y = 16'h200;
			16'h717f: y = 16'h200;
			16'h7180: y = 16'h200;
			16'h7181: y = 16'h200;
			16'h7182: y = 16'h200;
			16'h7183: y = 16'h200;
			16'h7184: y = 16'h200;
			16'h7185: y = 16'h200;
			16'h7186: y = 16'h200;
			16'h7187: y = 16'h200;
			16'h7188: y = 16'h200;
			16'h7189: y = 16'h200;
			16'h718a: y = 16'h200;
			16'h718b: y = 16'h200;
			16'h718c: y = 16'h200;
			16'h718d: y = 16'h200;
			16'h718e: y = 16'h200;
			16'h718f: y = 16'h200;
			16'h7190: y = 16'h200;
			16'h7191: y = 16'h200;
			16'h7192: y = 16'h200;
			16'h7193: y = 16'h200;
			16'h7194: y = 16'h200;
			16'h7195: y = 16'h200;
			16'h7196: y = 16'h200;
			16'h7197: y = 16'h200;
			16'h7198: y = 16'h200;
			16'h7199: y = 16'h200;
			16'h719a: y = 16'h200;
			16'h719b: y = 16'h200;
			16'h719c: y = 16'h200;
			16'h719d: y = 16'h200;
			16'h719e: y = 16'h200;
			16'h719f: y = 16'h200;
			16'h71a0: y = 16'h200;
			16'h71a1: y = 16'h200;
			16'h71a2: y = 16'h200;
			16'h71a3: y = 16'h200;
			16'h71a4: y = 16'h200;
			16'h71a5: y = 16'h200;
			16'h71a6: y = 16'h200;
			16'h71a7: y = 16'h200;
			16'h71a8: y = 16'h200;
			16'h71a9: y = 16'h200;
			16'h71aa: y = 16'h200;
			16'h71ab: y = 16'h200;
			16'h71ac: y = 16'h200;
			16'h71ad: y = 16'h200;
			16'h71ae: y = 16'h200;
			16'h71af: y = 16'h200;
			16'h71b0: y = 16'h200;
			16'h71b1: y = 16'h200;
			16'h71b2: y = 16'h200;
			16'h71b3: y = 16'h200;
			16'h71b4: y = 16'h200;
			16'h71b5: y = 16'h200;
			16'h71b6: y = 16'h200;
			16'h71b7: y = 16'h200;
			16'h71b8: y = 16'h200;
			16'h71b9: y = 16'h200;
			16'h71ba: y = 16'h200;
			16'h71bb: y = 16'h200;
			16'h71bc: y = 16'h200;
			16'h71bd: y = 16'h200;
			16'h71be: y = 16'h200;
			16'h71bf: y = 16'h200;
			16'h71c0: y = 16'h200;
			16'h71c1: y = 16'h200;
			16'h71c2: y = 16'h200;
			16'h71c3: y = 16'h200;
			16'h71c4: y = 16'h200;
			16'h71c5: y = 16'h200;
			16'h71c6: y = 16'h200;
			16'h71c7: y = 16'h200;
			16'h71c8: y = 16'h200;
			16'h71c9: y = 16'h200;
			16'h71ca: y = 16'h200;
			16'h71cb: y = 16'h200;
			16'h71cc: y = 16'h200;
			16'h71cd: y = 16'h200;
			16'h71ce: y = 16'h200;
			16'h71cf: y = 16'h200;
			16'h71d0: y = 16'h200;
			16'h71d1: y = 16'h200;
			16'h71d2: y = 16'h200;
			16'h71d3: y = 16'h200;
			16'h71d4: y = 16'h200;
			16'h71d5: y = 16'h200;
			16'h71d6: y = 16'h200;
			16'h71d7: y = 16'h200;
			16'h71d8: y = 16'h200;
			16'h71d9: y = 16'h200;
			16'h71da: y = 16'h200;
			16'h71db: y = 16'h200;
			16'h71dc: y = 16'h200;
			16'h71dd: y = 16'h200;
			16'h71de: y = 16'h200;
			16'h71df: y = 16'h200;
			16'h71e0: y = 16'h200;
			16'h71e1: y = 16'h200;
			16'h71e2: y = 16'h200;
			16'h71e3: y = 16'h200;
			16'h71e4: y = 16'h200;
			16'h71e5: y = 16'h200;
			16'h71e6: y = 16'h200;
			16'h71e7: y = 16'h200;
			16'h71e8: y = 16'h200;
			16'h71e9: y = 16'h200;
			16'h71ea: y = 16'h200;
			16'h71eb: y = 16'h200;
			16'h71ec: y = 16'h200;
			16'h71ed: y = 16'h200;
			16'h71ee: y = 16'h200;
			16'h71ef: y = 16'h200;
			16'h71f0: y = 16'h200;
			16'h71f1: y = 16'h200;
			16'h71f2: y = 16'h200;
			16'h71f3: y = 16'h200;
			16'h71f4: y = 16'h200;
			16'h71f5: y = 16'h200;
			16'h71f6: y = 16'h200;
			16'h71f7: y = 16'h200;
			16'h71f8: y = 16'h200;
			16'h71f9: y = 16'h200;
			16'h71fa: y = 16'h200;
			16'h71fb: y = 16'h200;
			16'h71fc: y = 16'h200;
			16'h71fd: y = 16'h200;
			16'h71fe: y = 16'h200;
			16'h71ff: y = 16'h200;
			16'h7200: y = 16'h200;
			16'h7201: y = 16'h200;
			16'h7202: y = 16'h200;
			16'h7203: y = 16'h200;
			16'h7204: y = 16'h200;
			16'h7205: y = 16'h200;
			16'h7206: y = 16'h200;
			16'h7207: y = 16'h200;
			16'h7208: y = 16'h200;
			16'h7209: y = 16'h200;
			16'h720a: y = 16'h200;
			16'h720b: y = 16'h200;
			16'h720c: y = 16'h200;
			16'h720d: y = 16'h200;
			16'h720e: y = 16'h200;
			16'h720f: y = 16'h200;
			16'h7210: y = 16'h200;
			16'h7211: y = 16'h200;
			16'h7212: y = 16'h200;
			16'h7213: y = 16'h200;
			16'h7214: y = 16'h200;
			16'h7215: y = 16'h200;
			16'h7216: y = 16'h200;
			16'h7217: y = 16'h200;
			16'h7218: y = 16'h200;
			16'h7219: y = 16'h200;
			16'h721a: y = 16'h200;
			16'h721b: y = 16'h200;
			16'h721c: y = 16'h200;
			16'h721d: y = 16'h200;
			16'h721e: y = 16'h200;
			16'h721f: y = 16'h200;
			16'h7220: y = 16'h200;
			16'h7221: y = 16'h200;
			16'h7222: y = 16'h200;
			16'h7223: y = 16'h200;
			16'h7224: y = 16'h200;
			16'h7225: y = 16'h200;
			16'h7226: y = 16'h200;
			16'h7227: y = 16'h200;
			16'h7228: y = 16'h200;
			16'h7229: y = 16'h200;
			16'h722a: y = 16'h200;
			16'h722b: y = 16'h200;
			16'h722c: y = 16'h200;
			16'h722d: y = 16'h200;
			16'h722e: y = 16'h200;
			16'h722f: y = 16'h200;
			16'h7230: y = 16'h200;
			16'h7231: y = 16'h200;
			16'h7232: y = 16'h200;
			16'h7233: y = 16'h200;
			16'h7234: y = 16'h200;
			16'h7235: y = 16'h200;
			16'h7236: y = 16'h200;
			16'h7237: y = 16'h200;
			16'h7238: y = 16'h200;
			16'h7239: y = 16'h200;
			16'h723a: y = 16'h200;
			16'h723b: y = 16'h200;
			16'h723c: y = 16'h200;
			16'h723d: y = 16'h200;
			16'h723e: y = 16'h200;
			16'h723f: y = 16'h200;
			16'h7240: y = 16'h200;
			16'h7241: y = 16'h200;
			16'h7242: y = 16'h200;
			16'h7243: y = 16'h200;
			16'h7244: y = 16'h200;
			16'h7245: y = 16'h200;
			16'h7246: y = 16'h200;
			16'h7247: y = 16'h200;
			16'h7248: y = 16'h200;
			16'h7249: y = 16'h200;
			16'h724a: y = 16'h200;
			16'h724b: y = 16'h200;
			16'h724c: y = 16'h200;
			16'h724d: y = 16'h200;
			16'h724e: y = 16'h200;
			16'h724f: y = 16'h200;
			16'h7250: y = 16'h200;
			16'h7251: y = 16'h200;
			16'h7252: y = 16'h200;
			16'h7253: y = 16'h200;
			16'h7254: y = 16'h200;
			16'h7255: y = 16'h200;
			16'h7256: y = 16'h200;
			16'h7257: y = 16'h200;
			16'h7258: y = 16'h200;
			16'h7259: y = 16'h200;
			16'h725a: y = 16'h200;
			16'h725b: y = 16'h200;
			16'h725c: y = 16'h200;
			16'h725d: y = 16'h200;
			16'h725e: y = 16'h200;
			16'h725f: y = 16'h200;
			16'h7260: y = 16'h200;
			16'h7261: y = 16'h200;
			16'h7262: y = 16'h200;
			16'h7263: y = 16'h200;
			16'h7264: y = 16'h200;
			16'h7265: y = 16'h200;
			16'h7266: y = 16'h200;
			16'h7267: y = 16'h200;
			16'h7268: y = 16'h200;
			16'h7269: y = 16'h200;
			16'h726a: y = 16'h200;
			16'h726b: y = 16'h200;
			16'h726c: y = 16'h200;
			16'h726d: y = 16'h200;
			16'h726e: y = 16'h200;
			16'h726f: y = 16'h200;
			16'h7270: y = 16'h200;
			16'h7271: y = 16'h200;
			16'h7272: y = 16'h200;
			16'h7273: y = 16'h200;
			16'h7274: y = 16'h200;
			16'h7275: y = 16'h200;
			16'h7276: y = 16'h200;
			16'h7277: y = 16'h200;
			16'h7278: y = 16'h200;
			16'h7279: y = 16'h200;
			16'h727a: y = 16'h200;
			16'h727b: y = 16'h200;
			16'h727c: y = 16'h200;
			16'h727d: y = 16'h200;
			16'h727e: y = 16'h200;
			16'h727f: y = 16'h200;
			16'h7280: y = 16'h200;
			16'h7281: y = 16'h200;
			16'h7282: y = 16'h200;
			16'h7283: y = 16'h200;
			16'h7284: y = 16'h200;
			16'h7285: y = 16'h200;
			16'h7286: y = 16'h200;
			16'h7287: y = 16'h200;
			16'h7288: y = 16'h200;
			16'h7289: y = 16'h200;
			16'h728a: y = 16'h200;
			16'h728b: y = 16'h200;
			16'h728c: y = 16'h200;
			16'h728d: y = 16'h200;
			16'h728e: y = 16'h200;
			16'h728f: y = 16'h200;
			16'h7290: y = 16'h200;
			16'h7291: y = 16'h200;
			16'h7292: y = 16'h200;
			16'h7293: y = 16'h200;
			16'h7294: y = 16'h200;
			16'h7295: y = 16'h200;
			16'h7296: y = 16'h200;
			16'h7297: y = 16'h200;
			16'h7298: y = 16'h200;
			16'h7299: y = 16'h200;
			16'h729a: y = 16'h200;
			16'h729b: y = 16'h200;
			16'h729c: y = 16'h200;
			16'h729d: y = 16'h200;
			16'h729e: y = 16'h200;
			16'h729f: y = 16'h200;
			16'h72a0: y = 16'h200;
			16'h72a1: y = 16'h200;
			16'h72a2: y = 16'h200;
			16'h72a3: y = 16'h200;
			16'h72a4: y = 16'h200;
			16'h72a5: y = 16'h200;
			16'h72a6: y = 16'h200;
			16'h72a7: y = 16'h200;
			16'h72a8: y = 16'h200;
			16'h72a9: y = 16'h200;
			16'h72aa: y = 16'h200;
			16'h72ab: y = 16'h200;
			16'h72ac: y = 16'h200;
			16'h72ad: y = 16'h200;
			16'h72ae: y = 16'h200;
			16'h72af: y = 16'h200;
			16'h72b0: y = 16'h200;
			16'h72b1: y = 16'h200;
			16'h72b2: y = 16'h200;
			16'h72b3: y = 16'h200;
			16'h72b4: y = 16'h200;
			16'h72b5: y = 16'h200;
			16'h72b6: y = 16'h200;
			16'h72b7: y = 16'h200;
			16'h72b8: y = 16'h200;
			16'h72b9: y = 16'h200;
			16'h72ba: y = 16'h200;
			16'h72bb: y = 16'h200;
			16'h72bc: y = 16'h200;
			16'h72bd: y = 16'h200;
			16'h72be: y = 16'h200;
			16'h72bf: y = 16'h200;
			16'h72c0: y = 16'h200;
			16'h72c1: y = 16'h200;
			16'h72c2: y = 16'h200;
			16'h72c3: y = 16'h200;
			16'h72c4: y = 16'h200;
			16'h72c5: y = 16'h200;
			16'h72c6: y = 16'h200;
			16'h72c7: y = 16'h200;
			16'h72c8: y = 16'h200;
			16'h72c9: y = 16'h200;
			16'h72ca: y = 16'h200;
			16'h72cb: y = 16'h200;
			16'h72cc: y = 16'h200;
			16'h72cd: y = 16'h200;
			16'h72ce: y = 16'h200;
			16'h72cf: y = 16'h200;
			16'h72d0: y = 16'h200;
			16'h72d1: y = 16'h200;
			16'h72d2: y = 16'h200;
			16'h72d3: y = 16'h200;
			16'h72d4: y = 16'h200;
			16'h72d5: y = 16'h200;
			16'h72d6: y = 16'h200;
			16'h72d7: y = 16'h200;
			16'h72d8: y = 16'h200;
			16'h72d9: y = 16'h200;
			16'h72da: y = 16'h200;
			16'h72db: y = 16'h200;
			16'h72dc: y = 16'h200;
			16'h72dd: y = 16'h200;
			16'h72de: y = 16'h200;
			16'h72df: y = 16'h200;
			16'h72e0: y = 16'h200;
			16'h72e1: y = 16'h200;
			16'h72e2: y = 16'h200;
			16'h72e3: y = 16'h200;
			16'h72e4: y = 16'h200;
			16'h72e5: y = 16'h200;
			16'h72e6: y = 16'h200;
			16'h72e7: y = 16'h200;
			16'h72e8: y = 16'h200;
			16'h72e9: y = 16'h200;
			16'h72ea: y = 16'h200;
			16'h72eb: y = 16'h200;
			16'h72ec: y = 16'h200;
			16'h72ed: y = 16'h200;
			16'h72ee: y = 16'h200;
			16'h72ef: y = 16'h200;
			16'h72f0: y = 16'h200;
			16'h72f1: y = 16'h200;
			16'h72f2: y = 16'h200;
			16'h72f3: y = 16'h200;
			16'h72f4: y = 16'h200;
			16'h72f5: y = 16'h200;
			16'h72f6: y = 16'h200;
			16'h72f7: y = 16'h200;
			16'h72f8: y = 16'h200;
			16'h72f9: y = 16'h200;
			16'h72fa: y = 16'h200;
			16'h72fb: y = 16'h200;
			16'h72fc: y = 16'h200;
			16'h72fd: y = 16'h200;
			16'h72fe: y = 16'h200;
			16'h72ff: y = 16'h200;
			16'h7300: y = 16'h200;
			16'h7301: y = 16'h200;
			16'h7302: y = 16'h200;
			16'h7303: y = 16'h200;
			16'h7304: y = 16'h200;
			16'h7305: y = 16'h200;
			16'h7306: y = 16'h200;
			16'h7307: y = 16'h200;
			16'h7308: y = 16'h200;
			16'h7309: y = 16'h200;
			16'h730a: y = 16'h200;
			16'h730b: y = 16'h200;
			16'h730c: y = 16'h200;
			16'h730d: y = 16'h200;
			16'h730e: y = 16'h200;
			16'h730f: y = 16'h200;
			16'h7310: y = 16'h200;
			16'h7311: y = 16'h200;
			16'h7312: y = 16'h200;
			16'h7313: y = 16'h200;
			16'h7314: y = 16'h200;
			16'h7315: y = 16'h200;
			16'h7316: y = 16'h200;
			16'h7317: y = 16'h200;
			16'h7318: y = 16'h200;
			16'h7319: y = 16'h200;
			16'h731a: y = 16'h200;
			16'h731b: y = 16'h200;
			16'h731c: y = 16'h200;
			16'h731d: y = 16'h200;
			16'h731e: y = 16'h200;
			16'h731f: y = 16'h200;
			16'h7320: y = 16'h200;
			16'h7321: y = 16'h200;
			16'h7322: y = 16'h200;
			16'h7323: y = 16'h200;
			16'h7324: y = 16'h200;
			16'h7325: y = 16'h200;
			16'h7326: y = 16'h200;
			16'h7327: y = 16'h200;
			16'h7328: y = 16'h200;
			16'h7329: y = 16'h200;
			16'h732a: y = 16'h200;
			16'h732b: y = 16'h200;
			16'h732c: y = 16'h200;
			16'h732d: y = 16'h200;
			16'h732e: y = 16'h200;
			16'h732f: y = 16'h200;
			16'h7330: y = 16'h200;
			16'h7331: y = 16'h200;
			16'h7332: y = 16'h200;
			16'h7333: y = 16'h200;
			16'h7334: y = 16'h200;
			16'h7335: y = 16'h200;
			16'h7336: y = 16'h200;
			16'h7337: y = 16'h200;
			16'h7338: y = 16'h200;
			16'h7339: y = 16'h200;
			16'h733a: y = 16'h200;
			16'h733b: y = 16'h200;
			16'h733c: y = 16'h200;
			16'h733d: y = 16'h200;
			16'h733e: y = 16'h200;
			16'h733f: y = 16'h200;
			16'h7340: y = 16'h200;
			16'h7341: y = 16'h200;
			16'h7342: y = 16'h200;
			16'h7343: y = 16'h200;
			16'h7344: y = 16'h200;
			16'h7345: y = 16'h200;
			16'h7346: y = 16'h200;
			16'h7347: y = 16'h200;
			16'h7348: y = 16'h200;
			16'h7349: y = 16'h200;
			16'h734a: y = 16'h200;
			16'h734b: y = 16'h200;
			16'h734c: y = 16'h200;
			16'h734d: y = 16'h200;
			16'h734e: y = 16'h200;
			16'h734f: y = 16'h200;
			16'h7350: y = 16'h200;
			16'h7351: y = 16'h200;
			16'h7352: y = 16'h200;
			16'h7353: y = 16'h200;
			16'h7354: y = 16'h200;
			16'h7355: y = 16'h200;
			16'h7356: y = 16'h200;
			16'h7357: y = 16'h200;
			16'h7358: y = 16'h200;
			16'h7359: y = 16'h200;
			16'h735a: y = 16'h200;
			16'h735b: y = 16'h200;
			16'h735c: y = 16'h200;
			16'h735d: y = 16'h200;
			16'h735e: y = 16'h200;
			16'h735f: y = 16'h200;
			16'h7360: y = 16'h200;
			16'h7361: y = 16'h200;
			16'h7362: y = 16'h200;
			16'h7363: y = 16'h200;
			16'h7364: y = 16'h200;
			16'h7365: y = 16'h200;
			16'h7366: y = 16'h200;
			16'h7367: y = 16'h200;
			16'h7368: y = 16'h200;
			16'h7369: y = 16'h200;
			16'h736a: y = 16'h200;
			16'h736b: y = 16'h200;
			16'h736c: y = 16'h200;
			16'h736d: y = 16'h200;
			16'h736e: y = 16'h200;
			16'h736f: y = 16'h200;
			16'h7370: y = 16'h200;
			16'h7371: y = 16'h200;
			16'h7372: y = 16'h200;
			16'h7373: y = 16'h200;
			16'h7374: y = 16'h200;
			16'h7375: y = 16'h200;
			16'h7376: y = 16'h200;
			16'h7377: y = 16'h200;
			16'h7378: y = 16'h200;
			16'h7379: y = 16'h200;
			16'h737a: y = 16'h200;
			16'h737b: y = 16'h200;
			16'h737c: y = 16'h200;
			16'h737d: y = 16'h200;
			16'h737e: y = 16'h200;
			16'h737f: y = 16'h200;
			16'h7380: y = 16'h200;
			16'h7381: y = 16'h200;
			16'h7382: y = 16'h200;
			16'h7383: y = 16'h200;
			16'h7384: y = 16'h200;
			16'h7385: y = 16'h200;
			16'h7386: y = 16'h200;
			16'h7387: y = 16'h200;
			16'h7388: y = 16'h200;
			16'h7389: y = 16'h200;
			16'h738a: y = 16'h200;
			16'h738b: y = 16'h200;
			16'h738c: y = 16'h200;
			16'h738d: y = 16'h200;
			16'h738e: y = 16'h200;
			16'h738f: y = 16'h200;
			16'h7390: y = 16'h200;
			16'h7391: y = 16'h200;
			16'h7392: y = 16'h200;
			16'h7393: y = 16'h200;
			16'h7394: y = 16'h200;
			16'h7395: y = 16'h200;
			16'h7396: y = 16'h200;
			16'h7397: y = 16'h200;
			16'h7398: y = 16'h200;
			16'h7399: y = 16'h200;
			16'h739a: y = 16'h200;
			16'h739b: y = 16'h200;
			16'h739c: y = 16'h200;
			16'h739d: y = 16'h200;
			16'h739e: y = 16'h200;
			16'h739f: y = 16'h200;
			16'h73a0: y = 16'h200;
			16'h73a1: y = 16'h200;
			16'h73a2: y = 16'h200;
			16'h73a3: y = 16'h200;
			16'h73a4: y = 16'h200;
			16'h73a5: y = 16'h200;
			16'h73a6: y = 16'h200;
			16'h73a7: y = 16'h200;
			16'h73a8: y = 16'h200;
			16'h73a9: y = 16'h200;
			16'h73aa: y = 16'h200;
			16'h73ab: y = 16'h200;
			16'h73ac: y = 16'h200;
			16'h73ad: y = 16'h200;
			16'h73ae: y = 16'h200;
			16'h73af: y = 16'h200;
			16'h73b0: y = 16'h200;
			16'h73b1: y = 16'h200;
			16'h73b2: y = 16'h200;
			16'h73b3: y = 16'h200;
			16'h73b4: y = 16'h200;
			16'h73b5: y = 16'h200;
			16'h73b6: y = 16'h200;
			16'h73b7: y = 16'h200;
			16'h73b8: y = 16'h200;
			16'h73b9: y = 16'h200;
			16'h73ba: y = 16'h200;
			16'h73bb: y = 16'h200;
			16'h73bc: y = 16'h200;
			16'h73bd: y = 16'h200;
			16'h73be: y = 16'h200;
			16'h73bf: y = 16'h200;
			16'h73c0: y = 16'h200;
			16'h73c1: y = 16'h200;
			16'h73c2: y = 16'h200;
			16'h73c3: y = 16'h200;
			16'h73c4: y = 16'h200;
			16'h73c5: y = 16'h200;
			16'h73c6: y = 16'h200;
			16'h73c7: y = 16'h200;
			16'h73c8: y = 16'h200;
			16'h73c9: y = 16'h200;
			16'h73ca: y = 16'h200;
			16'h73cb: y = 16'h200;
			16'h73cc: y = 16'h200;
			16'h73cd: y = 16'h200;
			16'h73ce: y = 16'h200;
			16'h73cf: y = 16'h200;
			16'h73d0: y = 16'h200;
			16'h73d1: y = 16'h200;
			16'h73d2: y = 16'h200;
			16'h73d3: y = 16'h200;
			16'h73d4: y = 16'h200;
			16'h73d5: y = 16'h200;
			16'h73d6: y = 16'h200;
			16'h73d7: y = 16'h200;
			16'h73d8: y = 16'h200;
			16'h73d9: y = 16'h200;
			16'h73da: y = 16'h200;
			16'h73db: y = 16'h200;
			16'h73dc: y = 16'h200;
			16'h73dd: y = 16'h200;
			16'h73de: y = 16'h200;
			16'h73df: y = 16'h200;
			16'h73e0: y = 16'h200;
			16'h73e1: y = 16'h200;
			16'h73e2: y = 16'h200;
			16'h73e3: y = 16'h200;
			16'h73e4: y = 16'h200;
			16'h73e5: y = 16'h200;
			16'h73e6: y = 16'h200;
			16'h73e7: y = 16'h200;
			16'h73e8: y = 16'h200;
			16'h73e9: y = 16'h200;
			16'h73ea: y = 16'h200;
			16'h73eb: y = 16'h200;
			16'h73ec: y = 16'h200;
			16'h73ed: y = 16'h200;
			16'h73ee: y = 16'h200;
			16'h73ef: y = 16'h200;
			16'h73f0: y = 16'h200;
			16'h73f1: y = 16'h200;
			16'h73f2: y = 16'h200;
			16'h73f3: y = 16'h200;
			16'h73f4: y = 16'h200;
			16'h73f5: y = 16'h200;
			16'h73f6: y = 16'h200;
			16'h73f7: y = 16'h200;
			16'h73f8: y = 16'h200;
			16'h73f9: y = 16'h200;
			16'h73fa: y = 16'h200;
			16'h73fb: y = 16'h200;
			16'h73fc: y = 16'h200;
			16'h73fd: y = 16'h200;
			16'h73fe: y = 16'h200;
			16'h73ff: y = 16'h200;
			16'h7400: y = 16'h200;
			16'h7401: y = 16'h200;
			16'h7402: y = 16'h200;
			16'h7403: y = 16'h200;
			16'h7404: y = 16'h200;
			16'h7405: y = 16'h200;
			16'h7406: y = 16'h200;
			16'h7407: y = 16'h200;
			16'h7408: y = 16'h200;
			16'h7409: y = 16'h200;
			16'h740a: y = 16'h200;
			16'h740b: y = 16'h200;
			16'h740c: y = 16'h200;
			16'h740d: y = 16'h200;
			16'h740e: y = 16'h200;
			16'h740f: y = 16'h200;
			16'h7410: y = 16'h200;
			16'h7411: y = 16'h200;
			16'h7412: y = 16'h200;
			16'h7413: y = 16'h200;
			16'h7414: y = 16'h200;
			16'h7415: y = 16'h200;
			16'h7416: y = 16'h200;
			16'h7417: y = 16'h200;
			16'h7418: y = 16'h200;
			16'h7419: y = 16'h200;
			16'h741a: y = 16'h200;
			16'h741b: y = 16'h200;
			16'h741c: y = 16'h200;
			16'h741d: y = 16'h200;
			16'h741e: y = 16'h200;
			16'h741f: y = 16'h200;
			16'h7420: y = 16'h200;
			16'h7421: y = 16'h200;
			16'h7422: y = 16'h200;
			16'h7423: y = 16'h200;
			16'h7424: y = 16'h200;
			16'h7425: y = 16'h200;
			16'h7426: y = 16'h200;
			16'h7427: y = 16'h200;
			16'h7428: y = 16'h200;
			16'h7429: y = 16'h200;
			16'h742a: y = 16'h200;
			16'h742b: y = 16'h200;
			16'h742c: y = 16'h200;
			16'h742d: y = 16'h200;
			16'h742e: y = 16'h200;
			16'h742f: y = 16'h200;
			16'h7430: y = 16'h200;
			16'h7431: y = 16'h200;
			16'h7432: y = 16'h200;
			16'h7433: y = 16'h200;
			16'h7434: y = 16'h200;
			16'h7435: y = 16'h200;
			16'h7436: y = 16'h200;
			16'h7437: y = 16'h200;
			16'h7438: y = 16'h200;
			16'h7439: y = 16'h200;
			16'h743a: y = 16'h200;
			16'h743b: y = 16'h200;
			16'h743c: y = 16'h200;
			16'h743d: y = 16'h200;
			16'h743e: y = 16'h200;
			16'h743f: y = 16'h200;
			16'h7440: y = 16'h200;
			16'h7441: y = 16'h200;
			16'h7442: y = 16'h200;
			16'h7443: y = 16'h200;
			16'h7444: y = 16'h200;
			16'h7445: y = 16'h200;
			16'h7446: y = 16'h200;
			16'h7447: y = 16'h200;
			16'h7448: y = 16'h200;
			16'h7449: y = 16'h200;
			16'h744a: y = 16'h200;
			16'h744b: y = 16'h200;
			16'h744c: y = 16'h200;
			16'h744d: y = 16'h200;
			16'h744e: y = 16'h200;
			16'h744f: y = 16'h200;
			16'h7450: y = 16'h200;
			16'h7451: y = 16'h200;
			16'h7452: y = 16'h200;
			16'h7453: y = 16'h200;
			16'h7454: y = 16'h200;
			16'h7455: y = 16'h200;
			16'h7456: y = 16'h200;
			16'h7457: y = 16'h200;
			16'h7458: y = 16'h200;
			16'h7459: y = 16'h200;
			16'h745a: y = 16'h200;
			16'h745b: y = 16'h200;
			16'h745c: y = 16'h200;
			16'h745d: y = 16'h200;
			16'h745e: y = 16'h200;
			16'h745f: y = 16'h200;
			16'h7460: y = 16'h200;
			16'h7461: y = 16'h200;
			16'h7462: y = 16'h200;
			16'h7463: y = 16'h200;
			16'h7464: y = 16'h200;
			16'h7465: y = 16'h200;
			16'h7466: y = 16'h200;
			16'h7467: y = 16'h200;
			16'h7468: y = 16'h200;
			16'h7469: y = 16'h200;
			16'h746a: y = 16'h200;
			16'h746b: y = 16'h200;
			16'h746c: y = 16'h200;
			16'h746d: y = 16'h200;
			16'h746e: y = 16'h200;
			16'h746f: y = 16'h200;
			16'h7470: y = 16'h200;
			16'h7471: y = 16'h200;
			16'h7472: y = 16'h200;
			16'h7473: y = 16'h200;
			16'h7474: y = 16'h200;
			16'h7475: y = 16'h200;
			16'h7476: y = 16'h200;
			16'h7477: y = 16'h200;
			16'h7478: y = 16'h200;
			16'h7479: y = 16'h200;
			16'h747a: y = 16'h200;
			16'h747b: y = 16'h200;
			16'h747c: y = 16'h200;
			16'h747d: y = 16'h200;
			16'h747e: y = 16'h200;
			16'h747f: y = 16'h200;
			16'h7480: y = 16'h200;
			16'h7481: y = 16'h200;
			16'h7482: y = 16'h200;
			16'h7483: y = 16'h200;
			16'h7484: y = 16'h200;
			16'h7485: y = 16'h200;
			16'h7486: y = 16'h200;
			16'h7487: y = 16'h200;
			16'h7488: y = 16'h200;
			16'h7489: y = 16'h200;
			16'h748a: y = 16'h200;
			16'h748b: y = 16'h200;
			16'h748c: y = 16'h200;
			16'h748d: y = 16'h200;
			16'h748e: y = 16'h200;
			16'h748f: y = 16'h200;
			16'h7490: y = 16'h200;
			16'h7491: y = 16'h200;
			16'h7492: y = 16'h200;
			16'h7493: y = 16'h200;
			16'h7494: y = 16'h200;
			16'h7495: y = 16'h200;
			16'h7496: y = 16'h200;
			16'h7497: y = 16'h200;
			16'h7498: y = 16'h200;
			16'h7499: y = 16'h200;
			16'h749a: y = 16'h200;
			16'h749b: y = 16'h200;
			16'h749c: y = 16'h200;
			16'h749d: y = 16'h200;
			16'h749e: y = 16'h200;
			16'h749f: y = 16'h200;
			16'h74a0: y = 16'h200;
			16'h74a1: y = 16'h200;
			16'h74a2: y = 16'h200;
			16'h74a3: y = 16'h200;
			16'h74a4: y = 16'h200;
			16'h74a5: y = 16'h200;
			16'h74a6: y = 16'h200;
			16'h74a7: y = 16'h200;
			16'h74a8: y = 16'h200;
			16'h74a9: y = 16'h200;
			16'h74aa: y = 16'h200;
			16'h74ab: y = 16'h200;
			16'h74ac: y = 16'h200;
			16'h74ad: y = 16'h200;
			16'h74ae: y = 16'h200;
			16'h74af: y = 16'h200;
			16'h74b0: y = 16'h200;
			16'h74b1: y = 16'h200;
			16'h74b2: y = 16'h200;
			16'h74b3: y = 16'h200;
			16'h74b4: y = 16'h200;
			16'h74b5: y = 16'h200;
			16'h74b6: y = 16'h200;
			16'h74b7: y = 16'h200;
			16'h74b8: y = 16'h200;
			16'h74b9: y = 16'h200;
			16'h74ba: y = 16'h200;
			16'h74bb: y = 16'h200;
			16'h74bc: y = 16'h200;
			16'h74bd: y = 16'h200;
			16'h74be: y = 16'h200;
			16'h74bf: y = 16'h200;
			16'h74c0: y = 16'h200;
			16'h74c1: y = 16'h200;
			16'h74c2: y = 16'h200;
			16'h74c3: y = 16'h200;
			16'h74c4: y = 16'h200;
			16'h74c5: y = 16'h200;
			16'h74c6: y = 16'h200;
			16'h74c7: y = 16'h200;
			16'h74c8: y = 16'h200;
			16'h74c9: y = 16'h200;
			16'h74ca: y = 16'h200;
			16'h74cb: y = 16'h200;
			16'h74cc: y = 16'h200;
			16'h74cd: y = 16'h200;
			16'h74ce: y = 16'h200;
			16'h74cf: y = 16'h200;
			16'h74d0: y = 16'h200;
			16'h74d1: y = 16'h200;
			16'h74d2: y = 16'h200;
			16'h74d3: y = 16'h200;
			16'h74d4: y = 16'h200;
			16'h74d5: y = 16'h200;
			16'h74d6: y = 16'h200;
			16'h74d7: y = 16'h200;
			16'h74d8: y = 16'h200;
			16'h74d9: y = 16'h200;
			16'h74da: y = 16'h200;
			16'h74db: y = 16'h200;
			16'h74dc: y = 16'h200;
			16'h74dd: y = 16'h200;
			16'h74de: y = 16'h200;
			16'h74df: y = 16'h200;
			16'h74e0: y = 16'h200;
			16'h74e1: y = 16'h200;
			16'h74e2: y = 16'h200;
			16'h74e3: y = 16'h200;
			16'h74e4: y = 16'h200;
			16'h74e5: y = 16'h200;
			16'h74e6: y = 16'h200;
			16'h74e7: y = 16'h200;
			16'h74e8: y = 16'h200;
			16'h74e9: y = 16'h200;
			16'h74ea: y = 16'h200;
			16'h74eb: y = 16'h200;
			16'h74ec: y = 16'h200;
			16'h74ed: y = 16'h200;
			16'h74ee: y = 16'h200;
			16'h74ef: y = 16'h200;
			16'h74f0: y = 16'h200;
			16'h74f1: y = 16'h200;
			16'h74f2: y = 16'h200;
			16'h74f3: y = 16'h200;
			16'h74f4: y = 16'h200;
			16'h74f5: y = 16'h200;
			16'h74f6: y = 16'h200;
			16'h74f7: y = 16'h200;
			16'h74f8: y = 16'h200;
			16'h74f9: y = 16'h200;
			16'h74fa: y = 16'h200;
			16'h74fb: y = 16'h200;
			16'h74fc: y = 16'h200;
			16'h74fd: y = 16'h200;
			16'h74fe: y = 16'h200;
			16'h74ff: y = 16'h200;
			16'h7500: y = 16'h200;
			16'h7501: y = 16'h200;
			16'h7502: y = 16'h200;
			16'h7503: y = 16'h200;
			16'h7504: y = 16'h200;
			16'h7505: y = 16'h200;
			16'h7506: y = 16'h200;
			16'h7507: y = 16'h200;
			16'h7508: y = 16'h200;
			16'h7509: y = 16'h200;
			16'h750a: y = 16'h200;
			16'h750b: y = 16'h200;
			16'h750c: y = 16'h200;
			16'h750d: y = 16'h200;
			16'h750e: y = 16'h200;
			16'h750f: y = 16'h200;
			16'h7510: y = 16'h200;
			16'h7511: y = 16'h200;
			16'h7512: y = 16'h200;
			16'h7513: y = 16'h200;
			16'h7514: y = 16'h200;
			16'h7515: y = 16'h200;
			16'h7516: y = 16'h200;
			16'h7517: y = 16'h200;
			16'h7518: y = 16'h200;
			16'h7519: y = 16'h200;
			16'h751a: y = 16'h200;
			16'h751b: y = 16'h200;
			16'h751c: y = 16'h200;
			16'h751d: y = 16'h200;
			16'h751e: y = 16'h200;
			16'h751f: y = 16'h200;
			16'h7520: y = 16'h200;
			16'h7521: y = 16'h200;
			16'h7522: y = 16'h200;
			16'h7523: y = 16'h200;
			16'h7524: y = 16'h200;
			16'h7525: y = 16'h200;
			16'h7526: y = 16'h200;
			16'h7527: y = 16'h200;
			16'h7528: y = 16'h200;
			16'h7529: y = 16'h200;
			16'h752a: y = 16'h200;
			16'h752b: y = 16'h200;
			16'h752c: y = 16'h200;
			16'h752d: y = 16'h200;
			16'h752e: y = 16'h200;
			16'h752f: y = 16'h200;
			16'h7530: y = 16'h200;
			16'h7531: y = 16'h200;
			16'h7532: y = 16'h200;
			16'h7533: y = 16'h200;
			16'h7534: y = 16'h200;
			16'h7535: y = 16'h200;
			16'h7536: y = 16'h200;
			16'h7537: y = 16'h200;
			16'h7538: y = 16'h200;
			16'h7539: y = 16'h200;
			16'h753a: y = 16'h200;
			16'h753b: y = 16'h200;
			16'h753c: y = 16'h200;
			16'h753d: y = 16'h200;
			16'h753e: y = 16'h200;
			16'h753f: y = 16'h200;
			16'h7540: y = 16'h200;
			16'h7541: y = 16'h200;
			16'h7542: y = 16'h200;
			16'h7543: y = 16'h200;
			16'h7544: y = 16'h200;
			16'h7545: y = 16'h200;
			16'h7546: y = 16'h200;
			16'h7547: y = 16'h200;
			16'h7548: y = 16'h200;
			16'h7549: y = 16'h200;
			16'h754a: y = 16'h200;
			16'h754b: y = 16'h200;
			16'h754c: y = 16'h200;
			16'h754d: y = 16'h200;
			16'h754e: y = 16'h200;
			16'h754f: y = 16'h200;
			16'h7550: y = 16'h200;
			16'h7551: y = 16'h200;
			16'h7552: y = 16'h200;
			16'h7553: y = 16'h200;
			16'h7554: y = 16'h200;
			16'h7555: y = 16'h200;
			16'h7556: y = 16'h200;
			16'h7557: y = 16'h200;
			16'h7558: y = 16'h200;
			16'h7559: y = 16'h200;
			16'h755a: y = 16'h200;
			16'h755b: y = 16'h200;
			16'h755c: y = 16'h200;
			16'h755d: y = 16'h200;
			16'h755e: y = 16'h200;
			16'h755f: y = 16'h200;
			16'h7560: y = 16'h200;
			16'h7561: y = 16'h200;
			16'h7562: y = 16'h200;
			16'h7563: y = 16'h200;
			16'h7564: y = 16'h200;
			16'h7565: y = 16'h200;
			16'h7566: y = 16'h200;
			16'h7567: y = 16'h200;
			16'h7568: y = 16'h200;
			16'h7569: y = 16'h200;
			16'h756a: y = 16'h200;
			16'h756b: y = 16'h200;
			16'h756c: y = 16'h200;
			16'h756d: y = 16'h200;
			16'h756e: y = 16'h200;
			16'h756f: y = 16'h200;
			16'h7570: y = 16'h200;
			16'h7571: y = 16'h200;
			16'h7572: y = 16'h200;
			16'h7573: y = 16'h200;
			16'h7574: y = 16'h200;
			16'h7575: y = 16'h200;
			16'h7576: y = 16'h200;
			16'h7577: y = 16'h200;
			16'h7578: y = 16'h200;
			16'h7579: y = 16'h200;
			16'h757a: y = 16'h200;
			16'h757b: y = 16'h200;
			16'h757c: y = 16'h200;
			16'h757d: y = 16'h200;
			16'h757e: y = 16'h200;
			16'h757f: y = 16'h200;
			16'h7580: y = 16'h200;
			16'h7581: y = 16'h200;
			16'h7582: y = 16'h200;
			16'h7583: y = 16'h200;
			16'h7584: y = 16'h200;
			16'h7585: y = 16'h200;
			16'h7586: y = 16'h200;
			16'h7587: y = 16'h200;
			16'h7588: y = 16'h200;
			16'h7589: y = 16'h200;
			16'h758a: y = 16'h200;
			16'h758b: y = 16'h200;
			16'h758c: y = 16'h200;
			16'h758d: y = 16'h200;
			16'h758e: y = 16'h200;
			16'h758f: y = 16'h200;
			16'h7590: y = 16'h200;
			16'h7591: y = 16'h200;
			16'h7592: y = 16'h200;
			16'h7593: y = 16'h200;
			16'h7594: y = 16'h200;
			16'h7595: y = 16'h200;
			16'h7596: y = 16'h200;
			16'h7597: y = 16'h200;
			16'h7598: y = 16'h200;
			16'h7599: y = 16'h200;
			16'h759a: y = 16'h200;
			16'h759b: y = 16'h200;
			16'h759c: y = 16'h200;
			16'h759d: y = 16'h200;
			16'h759e: y = 16'h200;
			16'h759f: y = 16'h200;
			16'h75a0: y = 16'h200;
			16'h75a1: y = 16'h200;
			16'h75a2: y = 16'h200;
			16'h75a3: y = 16'h200;
			16'h75a4: y = 16'h200;
			16'h75a5: y = 16'h200;
			16'h75a6: y = 16'h200;
			16'h75a7: y = 16'h200;
			16'h75a8: y = 16'h200;
			16'h75a9: y = 16'h200;
			16'h75aa: y = 16'h200;
			16'h75ab: y = 16'h200;
			16'h75ac: y = 16'h200;
			16'h75ad: y = 16'h200;
			16'h75ae: y = 16'h200;
			16'h75af: y = 16'h200;
			16'h75b0: y = 16'h200;
			16'h75b1: y = 16'h200;
			16'h75b2: y = 16'h200;
			16'h75b3: y = 16'h200;
			16'h75b4: y = 16'h200;
			16'h75b5: y = 16'h200;
			16'h75b6: y = 16'h200;
			16'h75b7: y = 16'h200;
			16'h75b8: y = 16'h200;
			16'h75b9: y = 16'h200;
			16'h75ba: y = 16'h200;
			16'h75bb: y = 16'h200;
			16'h75bc: y = 16'h200;
			16'h75bd: y = 16'h200;
			16'h75be: y = 16'h200;
			16'h75bf: y = 16'h200;
			16'h75c0: y = 16'h200;
			16'h75c1: y = 16'h200;
			16'h75c2: y = 16'h200;
			16'h75c3: y = 16'h200;
			16'h75c4: y = 16'h200;
			16'h75c5: y = 16'h200;
			16'h75c6: y = 16'h200;
			16'h75c7: y = 16'h200;
			16'h75c8: y = 16'h200;
			16'h75c9: y = 16'h200;
			16'h75ca: y = 16'h200;
			16'h75cb: y = 16'h200;
			16'h75cc: y = 16'h200;
			16'h75cd: y = 16'h200;
			16'h75ce: y = 16'h200;
			16'h75cf: y = 16'h200;
			16'h75d0: y = 16'h200;
			16'h75d1: y = 16'h200;
			16'h75d2: y = 16'h200;
			16'h75d3: y = 16'h200;
			16'h75d4: y = 16'h200;
			16'h75d5: y = 16'h200;
			16'h75d6: y = 16'h200;
			16'h75d7: y = 16'h200;
			16'h75d8: y = 16'h200;
			16'h75d9: y = 16'h200;
			16'h75da: y = 16'h200;
			16'h75db: y = 16'h200;
			16'h75dc: y = 16'h200;
			16'h75dd: y = 16'h200;
			16'h75de: y = 16'h200;
			16'h75df: y = 16'h200;
			16'h75e0: y = 16'h200;
			16'h75e1: y = 16'h200;
			16'h75e2: y = 16'h200;
			16'h75e3: y = 16'h200;
			16'h75e4: y = 16'h200;
			16'h75e5: y = 16'h200;
			16'h75e6: y = 16'h200;
			16'h75e7: y = 16'h200;
			16'h75e8: y = 16'h200;
			16'h75e9: y = 16'h200;
			16'h75ea: y = 16'h200;
			16'h75eb: y = 16'h200;
			16'h75ec: y = 16'h200;
			16'h75ed: y = 16'h200;
			16'h75ee: y = 16'h200;
			16'h75ef: y = 16'h200;
			16'h75f0: y = 16'h200;
			16'h75f1: y = 16'h200;
			16'h75f2: y = 16'h200;
			16'h75f3: y = 16'h200;
			16'h75f4: y = 16'h200;
			16'h75f5: y = 16'h200;
			16'h75f6: y = 16'h200;
			16'h75f7: y = 16'h200;
			16'h75f8: y = 16'h200;
			16'h75f9: y = 16'h200;
			16'h75fa: y = 16'h200;
			16'h75fb: y = 16'h200;
			16'h75fc: y = 16'h200;
			16'h75fd: y = 16'h200;
			16'h75fe: y = 16'h200;
			16'h75ff: y = 16'h200;
			16'h7600: y = 16'h200;
			16'h7601: y = 16'h200;
			16'h7602: y = 16'h200;
			16'h7603: y = 16'h200;
			16'h7604: y = 16'h200;
			16'h7605: y = 16'h200;
			16'h7606: y = 16'h200;
			16'h7607: y = 16'h200;
			16'h7608: y = 16'h200;
			16'h7609: y = 16'h200;
			16'h760a: y = 16'h200;
			16'h760b: y = 16'h200;
			16'h760c: y = 16'h200;
			16'h760d: y = 16'h200;
			16'h760e: y = 16'h200;
			16'h760f: y = 16'h200;
			16'h7610: y = 16'h200;
			16'h7611: y = 16'h200;
			16'h7612: y = 16'h200;
			16'h7613: y = 16'h200;
			16'h7614: y = 16'h200;
			16'h7615: y = 16'h200;
			16'h7616: y = 16'h200;
			16'h7617: y = 16'h200;
			16'h7618: y = 16'h200;
			16'h7619: y = 16'h200;
			16'h761a: y = 16'h200;
			16'h761b: y = 16'h200;
			16'h761c: y = 16'h200;
			16'h761d: y = 16'h200;
			16'h761e: y = 16'h200;
			16'h761f: y = 16'h200;
			16'h7620: y = 16'h200;
			16'h7621: y = 16'h200;
			16'h7622: y = 16'h200;
			16'h7623: y = 16'h200;
			16'h7624: y = 16'h200;
			16'h7625: y = 16'h200;
			16'h7626: y = 16'h200;
			16'h7627: y = 16'h200;
			16'h7628: y = 16'h200;
			16'h7629: y = 16'h200;
			16'h762a: y = 16'h200;
			16'h762b: y = 16'h200;
			16'h762c: y = 16'h200;
			16'h762d: y = 16'h200;
			16'h762e: y = 16'h200;
			16'h762f: y = 16'h200;
			16'h7630: y = 16'h200;
			16'h7631: y = 16'h200;
			16'h7632: y = 16'h200;
			16'h7633: y = 16'h200;
			16'h7634: y = 16'h200;
			16'h7635: y = 16'h200;
			16'h7636: y = 16'h200;
			16'h7637: y = 16'h200;
			16'h7638: y = 16'h200;
			16'h7639: y = 16'h200;
			16'h763a: y = 16'h200;
			16'h763b: y = 16'h200;
			16'h763c: y = 16'h200;
			16'h763d: y = 16'h200;
			16'h763e: y = 16'h200;
			16'h763f: y = 16'h200;
			16'h7640: y = 16'h200;
			16'h7641: y = 16'h200;
			16'h7642: y = 16'h200;
			16'h7643: y = 16'h200;
			16'h7644: y = 16'h200;
			16'h7645: y = 16'h200;
			16'h7646: y = 16'h200;
			16'h7647: y = 16'h200;
			16'h7648: y = 16'h200;
			16'h7649: y = 16'h200;
			16'h764a: y = 16'h200;
			16'h764b: y = 16'h200;
			16'h764c: y = 16'h200;
			16'h764d: y = 16'h200;
			16'h764e: y = 16'h200;
			16'h764f: y = 16'h200;
			16'h7650: y = 16'h200;
			16'h7651: y = 16'h200;
			16'h7652: y = 16'h200;
			16'h7653: y = 16'h200;
			16'h7654: y = 16'h200;
			16'h7655: y = 16'h200;
			16'h7656: y = 16'h200;
			16'h7657: y = 16'h200;
			16'h7658: y = 16'h200;
			16'h7659: y = 16'h200;
			16'h765a: y = 16'h200;
			16'h765b: y = 16'h200;
			16'h765c: y = 16'h200;
			16'h765d: y = 16'h200;
			16'h765e: y = 16'h200;
			16'h765f: y = 16'h200;
			16'h7660: y = 16'h200;
			16'h7661: y = 16'h200;
			16'h7662: y = 16'h200;
			16'h7663: y = 16'h200;
			16'h7664: y = 16'h200;
			16'h7665: y = 16'h200;
			16'h7666: y = 16'h200;
			16'h7667: y = 16'h200;
			16'h7668: y = 16'h200;
			16'h7669: y = 16'h200;
			16'h766a: y = 16'h200;
			16'h766b: y = 16'h200;
			16'h766c: y = 16'h200;
			16'h766d: y = 16'h200;
			16'h766e: y = 16'h200;
			16'h766f: y = 16'h200;
			16'h7670: y = 16'h200;
			16'h7671: y = 16'h200;
			16'h7672: y = 16'h200;
			16'h7673: y = 16'h200;
			16'h7674: y = 16'h200;
			16'h7675: y = 16'h200;
			16'h7676: y = 16'h200;
			16'h7677: y = 16'h200;
			16'h7678: y = 16'h200;
			16'h7679: y = 16'h200;
			16'h767a: y = 16'h200;
			16'h767b: y = 16'h200;
			16'h767c: y = 16'h200;
			16'h767d: y = 16'h200;
			16'h767e: y = 16'h200;
			16'h767f: y = 16'h200;
			16'h7680: y = 16'h200;
			16'h7681: y = 16'h200;
			16'h7682: y = 16'h200;
			16'h7683: y = 16'h200;
			16'h7684: y = 16'h200;
			16'h7685: y = 16'h200;
			16'h7686: y = 16'h200;
			16'h7687: y = 16'h200;
			16'h7688: y = 16'h200;
			16'h7689: y = 16'h200;
			16'h768a: y = 16'h200;
			16'h768b: y = 16'h200;
			16'h768c: y = 16'h200;
			16'h768d: y = 16'h200;
			16'h768e: y = 16'h200;
			16'h768f: y = 16'h200;
			16'h7690: y = 16'h200;
			16'h7691: y = 16'h200;
			16'h7692: y = 16'h200;
			16'h7693: y = 16'h200;
			16'h7694: y = 16'h200;
			16'h7695: y = 16'h200;
			16'h7696: y = 16'h200;
			16'h7697: y = 16'h200;
			16'h7698: y = 16'h200;
			16'h7699: y = 16'h200;
			16'h769a: y = 16'h200;
			16'h769b: y = 16'h200;
			16'h769c: y = 16'h200;
			16'h769d: y = 16'h200;
			16'h769e: y = 16'h200;
			16'h769f: y = 16'h200;
			16'h76a0: y = 16'h200;
			16'h76a1: y = 16'h200;
			16'h76a2: y = 16'h200;
			16'h76a3: y = 16'h200;
			16'h76a4: y = 16'h200;
			16'h76a5: y = 16'h200;
			16'h76a6: y = 16'h200;
			16'h76a7: y = 16'h200;
			16'h76a8: y = 16'h200;
			16'h76a9: y = 16'h200;
			16'h76aa: y = 16'h200;
			16'h76ab: y = 16'h200;
			16'h76ac: y = 16'h200;
			16'h76ad: y = 16'h200;
			16'h76ae: y = 16'h200;
			16'h76af: y = 16'h200;
			16'h76b0: y = 16'h200;
			16'h76b1: y = 16'h200;
			16'h76b2: y = 16'h200;
			16'h76b3: y = 16'h200;
			16'h76b4: y = 16'h200;
			16'h76b5: y = 16'h200;
			16'h76b6: y = 16'h200;
			16'h76b7: y = 16'h200;
			16'h76b8: y = 16'h200;
			16'h76b9: y = 16'h200;
			16'h76ba: y = 16'h200;
			16'h76bb: y = 16'h200;
			16'h76bc: y = 16'h200;
			16'h76bd: y = 16'h200;
			16'h76be: y = 16'h200;
			16'h76bf: y = 16'h200;
			16'h76c0: y = 16'h200;
			16'h76c1: y = 16'h200;
			16'h76c2: y = 16'h200;
			16'h76c3: y = 16'h200;
			16'h76c4: y = 16'h200;
			16'h76c5: y = 16'h200;
			16'h76c6: y = 16'h200;
			16'h76c7: y = 16'h200;
			16'h76c8: y = 16'h200;
			16'h76c9: y = 16'h200;
			16'h76ca: y = 16'h200;
			16'h76cb: y = 16'h200;
			16'h76cc: y = 16'h200;
			16'h76cd: y = 16'h200;
			16'h76ce: y = 16'h200;
			16'h76cf: y = 16'h200;
			16'h76d0: y = 16'h200;
			16'h76d1: y = 16'h200;
			16'h76d2: y = 16'h200;
			16'h76d3: y = 16'h200;
			16'h76d4: y = 16'h200;
			16'h76d5: y = 16'h200;
			16'h76d6: y = 16'h200;
			16'h76d7: y = 16'h200;
			16'h76d8: y = 16'h200;
			16'h76d9: y = 16'h200;
			16'h76da: y = 16'h200;
			16'h76db: y = 16'h200;
			16'h76dc: y = 16'h200;
			16'h76dd: y = 16'h200;
			16'h76de: y = 16'h200;
			16'h76df: y = 16'h200;
			16'h76e0: y = 16'h200;
			16'h76e1: y = 16'h200;
			16'h76e2: y = 16'h200;
			16'h76e3: y = 16'h200;
			16'h76e4: y = 16'h200;
			16'h76e5: y = 16'h200;
			16'h76e6: y = 16'h200;
			16'h76e7: y = 16'h200;
			16'h76e8: y = 16'h200;
			16'h76e9: y = 16'h200;
			16'h76ea: y = 16'h200;
			16'h76eb: y = 16'h200;
			16'h76ec: y = 16'h200;
			16'h76ed: y = 16'h200;
			16'h76ee: y = 16'h200;
			16'h76ef: y = 16'h200;
			16'h76f0: y = 16'h200;
			16'h76f1: y = 16'h200;
			16'h76f2: y = 16'h200;
			16'h76f3: y = 16'h200;
			16'h76f4: y = 16'h200;
			16'h76f5: y = 16'h200;
			16'h76f6: y = 16'h200;
			16'h76f7: y = 16'h200;
			16'h76f8: y = 16'h200;
			16'h76f9: y = 16'h200;
			16'h76fa: y = 16'h200;
			16'h76fb: y = 16'h200;
			16'h76fc: y = 16'h200;
			16'h76fd: y = 16'h200;
			16'h76fe: y = 16'h200;
			16'h76ff: y = 16'h200;
			16'h7700: y = 16'h200;
			16'h7701: y = 16'h200;
			16'h7702: y = 16'h200;
			16'h7703: y = 16'h200;
			16'h7704: y = 16'h200;
			16'h7705: y = 16'h200;
			16'h7706: y = 16'h200;
			16'h7707: y = 16'h200;
			16'h7708: y = 16'h200;
			16'h7709: y = 16'h200;
			16'h770a: y = 16'h200;
			16'h770b: y = 16'h200;
			16'h770c: y = 16'h200;
			16'h770d: y = 16'h200;
			16'h770e: y = 16'h200;
			16'h770f: y = 16'h200;
			16'h7710: y = 16'h200;
			16'h7711: y = 16'h200;
			16'h7712: y = 16'h200;
			16'h7713: y = 16'h200;
			16'h7714: y = 16'h200;
			16'h7715: y = 16'h200;
			16'h7716: y = 16'h200;
			16'h7717: y = 16'h200;
			16'h7718: y = 16'h200;
			16'h7719: y = 16'h200;
			16'h771a: y = 16'h200;
			16'h771b: y = 16'h200;
			16'h771c: y = 16'h200;
			16'h771d: y = 16'h200;
			16'h771e: y = 16'h200;
			16'h771f: y = 16'h200;
			16'h7720: y = 16'h200;
			16'h7721: y = 16'h200;
			16'h7722: y = 16'h200;
			16'h7723: y = 16'h200;
			16'h7724: y = 16'h200;
			16'h7725: y = 16'h200;
			16'h7726: y = 16'h200;
			16'h7727: y = 16'h200;
			16'h7728: y = 16'h200;
			16'h7729: y = 16'h200;
			16'h772a: y = 16'h200;
			16'h772b: y = 16'h200;
			16'h772c: y = 16'h200;
			16'h772d: y = 16'h200;
			16'h772e: y = 16'h200;
			16'h772f: y = 16'h200;
			16'h7730: y = 16'h200;
			16'h7731: y = 16'h200;
			16'h7732: y = 16'h200;
			16'h7733: y = 16'h200;
			16'h7734: y = 16'h200;
			16'h7735: y = 16'h200;
			16'h7736: y = 16'h200;
			16'h7737: y = 16'h200;
			16'h7738: y = 16'h200;
			16'h7739: y = 16'h200;
			16'h773a: y = 16'h200;
			16'h773b: y = 16'h200;
			16'h773c: y = 16'h200;
			16'h773d: y = 16'h200;
			16'h773e: y = 16'h200;
			16'h773f: y = 16'h200;
			16'h7740: y = 16'h200;
			16'h7741: y = 16'h200;
			16'h7742: y = 16'h200;
			16'h7743: y = 16'h200;
			16'h7744: y = 16'h200;
			16'h7745: y = 16'h200;
			16'h7746: y = 16'h200;
			16'h7747: y = 16'h200;
			16'h7748: y = 16'h200;
			16'h7749: y = 16'h200;
			16'h774a: y = 16'h200;
			16'h774b: y = 16'h200;
			16'h774c: y = 16'h200;
			16'h774d: y = 16'h200;
			16'h774e: y = 16'h200;
			16'h774f: y = 16'h200;
			16'h7750: y = 16'h200;
			16'h7751: y = 16'h200;
			16'h7752: y = 16'h200;
			16'h7753: y = 16'h200;
			16'h7754: y = 16'h200;
			16'h7755: y = 16'h200;
			16'h7756: y = 16'h200;
			16'h7757: y = 16'h200;
			16'h7758: y = 16'h200;
			16'h7759: y = 16'h200;
			16'h775a: y = 16'h200;
			16'h775b: y = 16'h200;
			16'h775c: y = 16'h200;
			16'h775d: y = 16'h200;
			16'h775e: y = 16'h200;
			16'h775f: y = 16'h200;
			16'h7760: y = 16'h200;
			16'h7761: y = 16'h200;
			16'h7762: y = 16'h200;
			16'h7763: y = 16'h200;
			16'h7764: y = 16'h200;
			16'h7765: y = 16'h200;
			16'h7766: y = 16'h200;
			16'h7767: y = 16'h200;
			16'h7768: y = 16'h200;
			16'h7769: y = 16'h200;
			16'h776a: y = 16'h200;
			16'h776b: y = 16'h200;
			16'h776c: y = 16'h200;
			16'h776d: y = 16'h200;
			16'h776e: y = 16'h200;
			16'h776f: y = 16'h200;
			16'h7770: y = 16'h200;
			16'h7771: y = 16'h200;
			16'h7772: y = 16'h200;
			16'h7773: y = 16'h200;
			16'h7774: y = 16'h200;
			16'h7775: y = 16'h200;
			16'h7776: y = 16'h200;
			16'h7777: y = 16'h200;
			16'h7778: y = 16'h200;
			16'h7779: y = 16'h200;
			16'h777a: y = 16'h200;
			16'h777b: y = 16'h200;
			16'h777c: y = 16'h200;
			16'h777d: y = 16'h200;
			16'h777e: y = 16'h200;
			16'h777f: y = 16'h200;
			16'h7780: y = 16'h200;
			16'h7781: y = 16'h200;
			16'h7782: y = 16'h200;
			16'h7783: y = 16'h200;
			16'h7784: y = 16'h200;
			16'h7785: y = 16'h200;
			16'h7786: y = 16'h200;
			16'h7787: y = 16'h200;
			16'h7788: y = 16'h200;
			16'h7789: y = 16'h200;
			16'h778a: y = 16'h200;
			16'h778b: y = 16'h200;
			16'h778c: y = 16'h200;
			16'h778d: y = 16'h200;
			16'h778e: y = 16'h200;
			16'h778f: y = 16'h200;
			16'h7790: y = 16'h200;
			16'h7791: y = 16'h200;
			16'h7792: y = 16'h200;
			16'h7793: y = 16'h200;
			16'h7794: y = 16'h200;
			16'h7795: y = 16'h200;
			16'h7796: y = 16'h200;
			16'h7797: y = 16'h200;
			16'h7798: y = 16'h200;
			16'h7799: y = 16'h200;
			16'h779a: y = 16'h200;
			16'h779b: y = 16'h200;
			16'h779c: y = 16'h200;
			16'h779d: y = 16'h200;
			16'h779e: y = 16'h200;
			16'h779f: y = 16'h200;
			16'h77a0: y = 16'h200;
			16'h77a1: y = 16'h200;
			16'h77a2: y = 16'h200;
			16'h77a3: y = 16'h200;
			16'h77a4: y = 16'h200;
			16'h77a5: y = 16'h200;
			16'h77a6: y = 16'h200;
			16'h77a7: y = 16'h200;
			16'h77a8: y = 16'h200;
			16'h77a9: y = 16'h200;
			16'h77aa: y = 16'h200;
			16'h77ab: y = 16'h200;
			16'h77ac: y = 16'h200;
			16'h77ad: y = 16'h200;
			16'h77ae: y = 16'h200;
			16'h77af: y = 16'h200;
			16'h77b0: y = 16'h200;
			16'h77b1: y = 16'h200;
			16'h77b2: y = 16'h200;
			16'h77b3: y = 16'h200;
			16'h77b4: y = 16'h200;
			16'h77b5: y = 16'h200;
			16'h77b6: y = 16'h200;
			16'h77b7: y = 16'h200;
			16'h77b8: y = 16'h200;
			16'h77b9: y = 16'h200;
			16'h77ba: y = 16'h200;
			16'h77bb: y = 16'h200;
			16'h77bc: y = 16'h200;
			16'h77bd: y = 16'h200;
			16'h77be: y = 16'h200;
			16'h77bf: y = 16'h200;
			16'h77c0: y = 16'h200;
			16'h77c1: y = 16'h200;
			16'h77c2: y = 16'h200;
			16'h77c3: y = 16'h200;
			16'h77c4: y = 16'h200;
			16'h77c5: y = 16'h200;
			16'h77c6: y = 16'h200;
			16'h77c7: y = 16'h200;
			16'h77c8: y = 16'h200;
			16'h77c9: y = 16'h200;
			16'h77ca: y = 16'h200;
			16'h77cb: y = 16'h200;
			16'h77cc: y = 16'h200;
			16'h77cd: y = 16'h200;
			16'h77ce: y = 16'h200;
			16'h77cf: y = 16'h200;
			16'h77d0: y = 16'h200;
			16'h77d1: y = 16'h200;
			16'h77d2: y = 16'h200;
			16'h77d3: y = 16'h200;
			16'h77d4: y = 16'h200;
			16'h77d5: y = 16'h200;
			16'h77d6: y = 16'h200;
			16'h77d7: y = 16'h200;
			16'h77d8: y = 16'h200;
			16'h77d9: y = 16'h200;
			16'h77da: y = 16'h200;
			16'h77db: y = 16'h200;
			16'h77dc: y = 16'h200;
			16'h77dd: y = 16'h200;
			16'h77de: y = 16'h200;
			16'h77df: y = 16'h200;
			16'h77e0: y = 16'h200;
			16'h77e1: y = 16'h200;
			16'h77e2: y = 16'h200;
			16'h77e3: y = 16'h200;
			16'h77e4: y = 16'h200;
			16'h77e5: y = 16'h200;
			16'h77e6: y = 16'h200;
			16'h77e7: y = 16'h200;
			16'h77e8: y = 16'h200;
			16'h77e9: y = 16'h200;
			16'h77ea: y = 16'h200;
			16'h77eb: y = 16'h200;
			16'h77ec: y = 16'h200;
			16'h77ed: y = 16'h200;
			16'h77ee: y = 16'h200;
			16'h77ef: y = 16'h200;
			16'h77f0: y = 16'h200;
			16'h77f1: y = 16'h200;
			16'h77f2: y = 16'h200;
			16'h77f3: y = 16'h200;
			16'h77f4: y = 16'h200;
			16'h77f5: y = 16'h200;
			16'h77f6: y = 16'h200;
			16'h77f7: y = 16'h200;
			16'h77f8: y = 16'h200;
			16'h77f9: y = 16'h200;
			16'h77fa: y = 16'h200;
			16'h77fb: y = 16'h200;
			16'h77fc: y = 16'h200;
			16'h77fd: y = 16'h200;
			16'h77fe: y = 16'h200;
			16'h77ff: y = 16'h200;
			16'h7800: y = 16'h200;
			16'h7801: y = 16'h200;
			16'h7802: y = 16'h200;
			16'h7803: y = 16'h200;
			16'h7804: y = 16'h200;
			16'h7805: y = 16'h200;
			16'h7806: y = 16'h200;
			16'h7807: y = 16'h200;
			16'h7808: y = 16'h200;
			16'h7809: y = 16'h200;
			16'h780a: y = 16'h200;
			16'h780b: y = 16'h200;
			16'h780c: y = 16'h200;
			16'h780d: y = 16'h200;
			16'h780e: y = 16'h200;
			16'h780f: y = 16'h200;
			16'h7810: y = 16'h200;
			16'h7811: y = 16'h200;
			16'h7812: y = 16'h200;
			16'h7813: y = 16'h200;
			16'h7814: y = 16'h200;
			16'h7815: y = 16'h200;
			16'h7816: y = 16'h200;
			16'h7817: y = 16'h200;
			16'h7818: y = 16'h200;
			16'h7819: y = 16'h200;
			16'h781a: y = 16'h200;
			16'h781b: y = 16'h200;
			16'h781c: y = 16'h200;
			16'h781d: y = 16'h200;
			16'h781e: y = 16'h200;
			16'h781f: y = 16'h200;
			16'h7820: y = 16'h200;
			16'h7821: y = 16'h200;
			16'h7822: y = 16'h200;
			16'h7823: y = 16'h200;
			16'h7824: y = 16'h200;
			16'h7825: y = 16'h200;
			16'h7826: y = 16'h200;
			16'h7827: y = 16'h200;
			16'h7828: y = 16'h200;
			16'h7829: y = 16'h200;
			16'h782a: y = 16'h200;
			16'h782b: y = 16'h200;
			16'h782c: y = 16'h200;
			16'h782d: y = 16'h200;
			16'h782e: y = 16'h200;
			16'h782f: y = 16'h200;
			16'h7830: y = 16'h200;
			16'h7831: y = 16'h200;
			16'h7832: y = 16'h200;
			16'h7833: y = 16'h200;
			16'h7834: y = 16'h200;
			16'h7835: y = 16'h200;
			16'h7836: y = 16'h200;
			16'h7837: y = 16'h200;
			16'h7838: y = 16'h200;
			16'h7839: y = 16'h200;
			16'h783a: y = 16'h200;
			16'h783b: y = 16'h200;
			16'h783c: y = 16'h200;
			16'h783d: y = 16'h200;
			16'h783e: y = 16'h200;
			16'h783f: y = 16'h200;
			16'h7840: y = 16'h200;
			16'h7841: y = 16'h200;
			16'h7842: y = 16'h200;
			16'h7843: y = 16'h200;
			16'h7844: y = 16'h200;
			16'h7845: y = 16'h200;
			16'h7846: y = 16'h200;
			16'h7847: y = 16'h200;
			16'h7848: y = 16'h200;
			16'h7849: y = 16'h200;
			16'h784a: y = 16'h200;
			16'h784b: y = 16'h200;
			16'h784c: y = 16'h200;
			16'h784d: y = 16'h200;
			16'h784e: y = 16'h200;
			16'h784f: y = 16'h200;
			16'h7850: y = 16'h200;
			16'h7851: y = 16'h200;
			16'h7852: y = 16'h200;
			16'h7853: y = 16'h200;
			16'h7854: y = 16'h200;
			16'h7855: y = 16'h200;
			16'h7856: y = 16'h200;
			16'h7857: y = 16'h200;
			16'h7858: y = 16'h200;
			16'h7859: y = 16'h200;
			16'h785a: y = 16'h200;
			16'h785b: y = 16'h200;
			16'h785c: y = 16'h200;
			16'h785d: y = 16'h200;
			16'h785e: y = 16'h200;
			16'h785f: y = 16'h200;
			16'h7860: y = 16'h200;
			16'h7861: y = 16'h200;
			16'h7862: y = 16'h200;
			16'h7863: y = 16'h200;
			16'h7864: y = 16'h200;
			16'h7865: y = 16'h200;
			16'h7866: y = 16'h200;
			16'h7867: y = 16'h200;
			16'h7868: y = 16'h200;
			16'h7869: y = 16'h200;
			16'h786a: y = 16'h200;
			16'h786b: y = 16'h200;
			16'h786c: y = 16'h200;
			16'h786d: y = 16'h200;
			16'h786e: y = 16'h200;
			16'h786f: y = 16'h200;
			16'h7870: y = 16'h200;
			16'h7871: y = 16'h200;
			16'h7872: y = 16'h200;
			16'h7873: y = 16'h200;
			16'h7874: y = 16'h200;
			16'h7875: y = 16'h200;
			16'h7876: y = 16'h200;
			16'h7877: y = 16'h200;
			16'h7878: y = 16'h200;
			16'h7879: y = 16'h200;
			16'h787a: y = 16'h200;
			16'h787b: y = 16'h200;
			16'h787c: y = 16'h200;
			16'h787d: y = 16'h200;
			16'h787e: y = 16'h200;
			16'h787f: y = 16'h200;
			16'h7880: y = 16'h200;
			16'h7881: y = 16'h200;
			16'h7882: y = 16'h200;
			16'h7883: y = 16'h200;
			16'h7884: y = 16'h200;
			16'h7885: y = 16'h200;
			16'h7886: y = 16'h200;
			16'h7887: y = 16'h200;
			16'h7888: y = 16'h200;
			16'h7889: y = 16'h200;
			16'h788a: y = 16'h200;
			16'h788b: y = 16'h200;
			16'h788c: y = 16'h200;
			16'h788d: y = 16'h200;
			16'h788e: y = 16'h200;
			16'h788f: y = 16'h200;
			16'h7890: y = 16'h200;
			16'h7891: y = 16'h200;
			16'h7892: y = 16'h200;
			16'h7893: y = 16'h200;
			16'h7894: y = 16'h200;
			16'h7895: y = 16'h200;
			16'h7896: y = 16'h200;
			16'h7897: y = 16'h200;
			16'h7898: y = 16'h200;
			16'h7899: y = 16'h200;
			16'h789a: y = 16'h200;
			16'h789b: y = 16'h200;
			16'h789c: y = 16'h200;
			16'h789d: y = 16'h200;
			16'h789e: y = 16'h200;
			16'h789f: y = 16'h200;
			16'h78a0: y = 16'h200;
			16'h78a1: y = 16'h200;
			16'h78a2: y = 16'h200;
			16'h78a3: y = 16'h200;
			16'h78a4: y = 16'h200;
			16'h78a5: y = 16'h200;
			16'h78a6: y = 16'h200;
			16'h78a7: y = 16'h200;
			16'h78a8: y = 16'h200;
			16'h78a9: y = 16'h200;
			16'h78aa: y = 16'h200;
			16'h78ab: y = 16'h200;
			16'h78ac: y = 16'h200;
			16'h78ad: y = 16'h200;
			16'h78ae: y = 16'h200;
			16'h78af: y = 16'h200;
			16'h78b0: y = 16'h200;
			16'h78b1: y = 16'h200;
			16'h78b2: y = 16'h200;
			16'h78b3: y = 16'h200;
			16'h78b4: y = 16'h200;
			16'h78b5: y = 16'h200;
			16'h78b6: y = 16'h200;
			16'h78b7: y = 16'h200;
			16'h78b8: y = 16'h200;
			16'h78b9: y = 16'h200;
			16'h78ba: y = 16'h200;
			16'h78bb: y = 16'h200;
			16'h78bc: y = 16'h200;
			16'h78bd: y = 16'h200;
			16'h78be: y = 16'h200;
			16'h78bf: y = 16'h200;
			16'h78c0: y = 16'h200;
			16'h78c1: y = 16'h200;
			16'h78c2: y = 16'h200;
			16'h78c3: y = 16'h200;
			16'h78c4: y = 16'h200;
			16'h78c5: y = 16'h200;
			16'h78c6: y = 16'h200;
			16'h78c7: y = 16'h200;
			16'h78c8: y = 16'h200;
			16'h78c9: y = 16'h200;
			16'h78ca: y = 16'h200;
			16'h78cb: y = 16'h200;
			16'h78cc: y = 16'h200;
			16'h78cd: y = 16'h200;
			16'h78ce: y = 16'h200;
			16'h78cf: y = 16'h200;
			16'h78d0: y = 16'h200;
			16'h78d1: y = 16'h200;
			16'h78d2: y = 16'h200;
			16'h78d3: y = 16'h200;
			16'h78d4: y = 16'h200;
			16'h78d5: y = 16'h200;
			16'h78d6: y = 16'h200;
			16'h78d7: y = 16'h200;
			16'h78d8: y = 16'h200;
			16'h78d9: y = 16'h200;
			16'h78da: y = 16'h200;
			16'h78db: y = 16'h200;
			16'h78dc: y = 16'h200;
			16'h78dd: y = 16'h200;
			16'h78de: y = 16'h200;
			16'h78df: y = 16'h200;
			16'h78e0: y = 16'h200;
			16'h78e1: y = 16'h200;
			16'h78e2: y = 16'h200;
			16'h78e3: y = 16'h200;
			16'h78e4: y = 16'h200;
			16'h78e5: y = 16'h200;
			16'h78e6: y = 16'h200;
			16'h78e7: y = 16'h200;
			16'h78e8: y = 16'h200;
			16'h78e9: y = 16'h200;
			16'h78ea: y = 16'h200;
			16'h78eb: y = 16'h200;
			16'h78ec: y = 16'h200;
			16'h78ed: y = 16'h200;
			16'h78ee: y = 16'h200;
			16'h78ef: y = 16'h200;
			16'h78f0: y = 16'h200;
			16'h78f1: y = 16'h200;
			16'h78f2: y = 16'h200;
			16'h78f3: y = 16'h200;
			16'h78f4: y = 16'h200;
			16'h78f5: y = 16'h200;
			16'h78f6: y = 16'h200;
			16'h78f7: y = 16'h200;
			16'h78f8: y = 16'h200;
			16'h78f9: y = 16'h200;
			16'h78fa: y = 16'h200;
			16'h78fb: y = 16'h200;
			16'h78fc: y = 16'h200;
			16'h78fd: y = 16'h200;
			16'h78fe: y = 16'h200;
			16'h78ff: y = 16'h200;
			16'h7900: y = 16'h200;
			16'h7901: y = 16'h200;
			16'h7902: y = 16'h200;
			16'h7903: y = 16'h200;
			16'h7904: y = 16'h200;
			16'h7905: y = 16'h200;
			16'h7906: y = 16'h200;
			16'h7907: y = 16'h200;
			16'h7908: y = 16'h200;
			16'h7909: y = 16'h200;
			16'h790a: y = 16'h200;
			16'h790b: y = 16'h200;
			16'h790c: y = 16'h200;
			16'h790d: y = 16'h200;
			16'h790e: y = 16'h200;
			16'h790f: y = 16'h200;
			16'h7910: y = 16'h200;
			16'h7911: y = 16'h200;
			16'h7912: y = 16'h200;
			16'h7913: y = 16'h200;
			16'h7914: y = 16'h200;
			16'h7915: y = 16'h200;
			16'h7916: y = 16'h200;
			16'h7917: y = 16'h200;
			16'h7918: y = 16'h200;
			16'h7919: y = 16'h200;
			16'h791a: y = 16'h200;
			16'h791b: y = 16'h200;
			16'h791c: y = 16'h200;
			16'h791d: y = 16'h200;
			16'h791e: y = 16'h200;
			16'h791f: y = 16'h200;
			16'h7920: y = 16'h200;
			16'h7921: y = 16'h200;
			16'h7922: y = 16'h200;
			16'h7923: y = 16'h200;
			16'h7924: y = 16'h200;
			16'h7925: y = 16'h200;
			16'h7926: y = 16'h200;
			16'h7927: y = 16'h200;
			16'h7928: y = 16'h200;
			16'h7929: y = 16'h200;
			16'h792a: y = 16'h200;
			16'h792b: y = 16'h200;
			16'h792c: y = 16'h200;
			16'h792d: y = 16'h200;
			16'h792e: y = 16'h200;
			16'h792f: y = 16'h200;
			16'h7930: y = 16'h200;
			16'h7931: y = 16'h200;
			16'h7932: y = 16'h200;
			16'h7933: y = 16'h200;
			16'h7934: y = 16'h200;
			16'h7935: y = 16'h200;
			16'h7936: y = 16'h200;
			16'h7937: y = 16'h200;
			16'h7938: y = 16'h200;
			16'h7939: y = 16'h200;
			16'h793a: y = 16'h200;
			16'h793b: y = 16'h200;
			16'h793c: y = 16'h200;
			16'h793d: y = 16'h200;
			16'h793e: y = 16'h200;
			16'h793f: y = 16'h200;
			16'h7940: y = 16'h200;
			16'h7941: y = 16'h200;
			16'h7942: y = 16'h200;
			16'h7943: y = 16'h200;
			16'h7944: y = 16'h200;
			16'h7945: y = 16'h200;
			16'h7946: y = 16'h200;
			16'h7947: y = 16'h200;
			16'h7948: y = 16'h200;
			16'h7949: y = 16'h200;
			16'h794a: y = 16'h200;
			16'h794b: y = 16'h200;
			16'h794c: y = 16'h200;
			16'h794d: y = 16'h200;
			16'h794e: y = 16'h200;
			16'h794f: y = 16'h200;
			16'h7950: y = 16'h200;
			16'h7951: y = 16'h200;
			16'h7952: y = 16'h200;
			16'h7953: y = 16'h200;
			16'h7954: y = 16'h200;
			16'h7955: y = 16'h200;
			16'h7956: y = 16'h200;
			16'h7957: y = 16'h200;
			16'h7958: y = 16'h200;
			16'h7959: y = 16'h200;
			16'h795a: y = 16'h200;
			16'h795b: y = 16'h200;
			16'h795c: y = 16'h200;
			16'h795d: y = 16'h200;
			16'h795e: y = 16'h200;
			16'h795f: y = 16'h200;
			16'h7960: y = 16'h200;
			16'h7961: y = 16'h200;
			16'h7962: y = 16'h200;
			16'h7963: y = 16'h200;
			16'h7964: y = 16'h200;
			16'h7965: y = 16'h200;
			16'h7966: y = 16'h200;
			16'h7967: y = 16'h200;
			16'h7968: y = 16'h200;
			16'h7969: y = 16'h200;
			16'h796a: y = 16'h200;
			16'h796b: y = 16'h200;
			16'h796c: y = 16'h200;
			16'h796d: y = 16'h200;
			16'h796e: y = 16'h200;
			16'h796f: y = 16'h200;
			16'h7970: y = 16'h200;
			16'h7971: y = 16'h200;
			16'h7972: y = 16'h200;
			16'h7973: y = 16'h200;
			16'h7974: y = 16'h200;
			16'h7975: y = 16'h200;
			16'h7976: y = 16'h200;
			16'h7977: y = 16'h200;
			16'h7978: y = 16'h200;
			16'h7979: y = 16'h200;
			16'h797a: y = 16'h200;
			16'h797b: y = 16'h200;
			16'h797c: y = 16'h200;
			16'h797d: y = 16'h200;
			16'h797e: y = 16'h200;
			16'h797f: y = 16'h200;
			16'h7980: y = 16'h200;
			16'h7981: y = 16'h200;
			16'h7982: y = 16'h200;
			16'h7983: y = 16'h200;
			16'h7984: y = 16'h200;
			16'h7985: y = 16'h200;
			16'h7986: y = 16'h200;
			16'h7987: y = 16'h200;
			16'h7988: y = 16'h200;
			16'h7989: y = 16'h200;
			16'h798a: y = 16'h200;
			16'h798b: y = 16'h200;
			16'h798c: y = 16'h200;
			16'h798d: y = 16'h200;
			16'h798e: y = 16'h200;
			16'h798f: y = 16'h200;
			16'h7990: y = 16'h200;
			16'h7991: y = 16'h200;
			16'h7992: y = 16'h200;
			16'h7993: y = 16'h200;
			16'h7994: y = 16'h200;
			16'h7995: y = 16'h200;
			16'h7996: y = 16'h200;
			16'h7997: y = 16'h200;
			16'h7998: y = 16'h200;
			16'h7999: y = 16'h200;
			16'h799a: y = 16'h200;
			16'h799b: y = 16'h200;
			16'h799c: y = 16'h200;
			16'h799d: y = 16'h200;
			16'h799e: y = 16'h200;
			16'h799f: y = 16'h200;
			16'h79a0: y = 16'h200;
			16'h79a1: y = 16'h200;
			16'h79a2: y = 16'h200;
			16'h79a3: y = 16'h200;
			16'h79a4: y = 16'h200;
			16'h79a5: y = 16'h200;
			16'h79a6: y = 16'h200;
			16'h79a7: y = 16'h200;
			16'h79a8: y = 16'h200;
			16'h79a9: y = 16'h200;
			16'h79aa: y = 16'h200;
			16'h79ab: y = 16'h200;
			16'h79ac: y = 16'h200;
			16'h79ad: y = 16'h200;
			16'h79ae: y = 16'h200;
			16'h79af: y = 16'h200;
			16'h79b0: y = 16'h200;
			16'h79b1: y = 16'h200;
			16'h79b2: y = 16'h200;
			16'h79b3: y = 16'h200;
			16'h79b4: y = 16'h200;
			16'h79b5: y = 16'h200;
			16'h79b6: y = 16'h200;
			16'h79b7: y = 16'h200;
			16'h79b8: y = 16'h200;
			16'h79b9: y = 16'h200;
			16'h79ba: y = 16'h200;
			16'h79bb: y = 16'h200;
			16'h79bc: y = 16'h200;
			16'h79bd: y = 16'h200;
			16'h79be: y = 16'h200;
			16'h79bf: y = 16'h200;
			16'h79c0: y = 16'h200;
			16'h79c1: y = 16'h200;
			16'h79c2: y = 16'h200;
			16'h79c3: y = 16'h200;
			16'h79c4: y = 16'h200;
			16'h79c5: y = 16'h200;
			16'h79c6: y = 16'h200;
			16'h79c7: y = 16'h200;
			16'h79c8: y = 16'h200;
			16'h79c9: y = 16'h200;
			16'h79ca: y = 16'h200;
			16'h79cb: y = 16'h200;
			16'h79cc: y = 16'h200;
			16'h79cd: y = 16'h200;
			16'h79ce: y = 16'h200;
			16'h79cf: y = 16'h200;
			16'h79d0: y = 16'h200;
			16'h79d1: y = 16'h200;
			16'h79d2: y = 16'h200;
			16'h79d3: y = 16'h200;
			16'h79d4: y = 16'h200;
			16'h79d5: y = 16'h200;
			16'h79d6: y = 16'h200;
			16'h79d7: y = 16'h200;
			16'h79d8: y = 16'h200;
			16'h79d9: y = 16'h200;
			16'h79da: y = 16'h200;
			16'h79db: y = 16'h200;
			16'h79dc: y = 16'h200;
			16'h79dd: y = 16'h200;
			16'h79de: y = 16'h200;
			16'h79df: y = 16'h200;
			16'h79e0: y = 16'h200;
			16'h79e1: y = 16'h200;
			16'h79e2: y = 16'h200;
			16'h79e3: y = 16'h200;
			16'h79e4: y = 16'h200;
			16'h79e5: y = 16'h200;
			16'h79e6: y = 16'h200;
			16'h79e7: y = 16'h200;
			16'h79e8: y = 16'h200;
			16'h79e9: y = 16'h200;
			16'h79ea: y = 16'h200;
			16'h79eb: y = 16'h200;
			16'h79ec: y = 16'h200;
			16'h79ed: y = 16'h200;
			16'h79ee: y = 16'h200;
			16'h79ef: y = 16'h200;
			16'h79f0: y = 16'h200;
			16'h79f1: y = 16'h200;
			16'h79f2: y = 16'h200;
			16'h79f3: y = 16'h200;
			16'h79f4: y = 16'h200;
			16'h79f5: y = 16'h200;
			16'h79f6: y = 16'h200;
			16'h79f7: y = 16'h200;
			16'h79f8: y = 16'h200;
			16'h79f9: y = 16'h200;
			16'h79fa: y = 16'h200;
			16'h79fb: y = 16'h200;
			16'h79fc: y = 16'h200;
			16'h79fd: y = 16'h200;
			16'h79fe: y = 16'h200;
			16'h79ff: y = 16'h200;
			16'h7a00: y = 16'h200;
			16'h7a01: y = 16'h200;
			16'h7a02: y = 16'h200;
			16'h7a03: y = 16'h200;
			16'h7a04: y = 16'h200;
			16'h7a05: y = 16'h200;
			16'h7a06: y = 16'h200;
			16'h7a07: y = 16'h200;
			16'h7a08: y = 16'h200;
			16'h7a09: y = 16'h200;
			16'h7a0a: y = 16'h200;
			16'h7a0b: y = 16'h200;
			16'h7a0c: y = 16'h200;
			16'h7a0d: y = 16'h200;
			16'h7a0e: y = 16'h200;
			16'h7a0f: y = 16'h200;
			16'h7a10: y = 16'h200;
			16'h7a11: y = 16'h200;
			16'h7a12: y = 16'h200;
			16'h7a13: y = 16'h200;
			16'h7a14: y = 16'h200;
			16'h7a15: y = 16'h200;
			16'h7a16: y = 16'h200;
			16'h7a17: y = 16'h200;
			16'h7a18: y = 16'h200;
			16'h7a19: y = 16'h200;
			16'h7a1a: y = 16'h200;
			16'h7a1b: y = 16'h200;
			16'h7a1c: y = 16'h200;
			16'h7a1d: y = 16'h200;
			16'h7a1e: y = 16'h200;
			16'h7a1f: y = 16'h200;
			16'h7a20: y = 16'h200;
			16'h7a21: y = 16'h200;
			16'h7a22: y = 16'h200;
			16'h7a23: y = 16'h200;
			16'h7a24: y = 16'h200;
			16'h7a25: y = 16'h200;
			16'h7a26: y = 16'h200;
			16'h7a27: y = 16'h200;
			16'h7a28: y = 16'h200;
			16'h7a29: y = 16'h200;
			16'h7a2a: y = 16'h200;
			16'h7a2b: y = 16'h200;
			16'h7a2c: y = 16'h200;
			16'h7a2d: y = 16'h200;
			16'h7a2e: y = 16'h200;
			16'h7a2f: y = 16'h200;
			16'h7a30: y = 16'h200;
			16'h7a31: y = 16'h200;
			16'h7a32: y = 16'h200;
			16'h7a33: y = 16'h200;
			16'h7a34: y = 16'h200;
			16'h7a35: y = 16'h200;
			16'h7a36: y = 16'h200;
			16'h7a37: y = 16'h200;
			16'h7a38: y = 16'h200;
			16'h7a39: y = 16'h200;
			16'h7a3a: y = 16'h200;
			16'h7a3b: y = 16'h200;
			16'h7a3c: y = 16'h200;
			16'h7a3d: y = 16'h200;
			16'h7a3e: y = 16'h200;
			16'h7a3f: y = 16'h200;
			16'h7a40: y = 16'h200;
			16'h7a41: y = 16'h200;
			16'h7a42: y = 16'h200;
			16'h7a43: y = 16'h200;
			16'h7a44: y = 16'h200;
			16'h7a45: y = 16'h200;
			16'h7a46: y = 16'h200;
			16'h7a47: y = 16'h200;
			16'h7a48: y = 16'h200;
			16'h7a49: y = 16'h200;
			16'h7a4a: y = 16'h200;
			16'h7a4b: y = 16'h200;
			16'h7a4c: y = 16'h200;
			16'h7a4d: y = 16'h200;
			16'h7a4e: y = 16'h200;
			16'h7a4f: y = 16'h200;
			16'h7a50: y = 16'h200;
			16'h7a51: y = 16'h200;
			16'h7a52: y = 16'h200;
			16'h7a53: y = 16'h200;
			16'h7a54: y = 16'h200;
			16'h7a55: y = 16'h200;
			16'h7a56: y = 16'h200;
			16'h7a57: y = 16'h200;
			16'h7a58: y = 16'h200;
			16'h7a59: y = 16'h200;
			16'h7a5a: y = 16'h200;
			16'h7a5b: y = 16'h200;
			16'h7a5c: y = 16'h200;
			16'h7a5d: y = 16'h200;
			16'h7a5e: y = 16'h200;
			16'h7a5f: y = 16'h200;
			16'h7a60: y = 16'h200;
			16'h7a61: y = 16'h200;
			16'h7a62: y = 16'h200;
			16'h7a63: y = 16'h200;
			16'h7a64: y = 16'h200;
			16'h7a65: y = 16'h200;
			16'h7a66: y = 16'h200;
			16'h7a67: y = 16'h200;
			16'h7a68: y = 16'h200;
			16'h7a69: y = 16'h200;
			16'h7a6a: y = 16'h200;
			16'h7a6b: y = 16'h200;
			16'h7a6c: y = 16'h200;
			16'h7a6d: y = 16'h200;
			16'h7a6e: y = 16'h200;
			16'h7a6f: y = 16'h200;
			16'h7a70: y = 16'h200;
			16'h7a71: y = 16'h200;
			16'h7a72: y = 16'h200;
			16'h7a73: y = 16'h200;
			16'h7a74: y = 16'h200;
			16'h7a75: y = 16'h200;
			16'h7a76: y = 16'h200;
			16'h7a77: y = 16'h200;
			16'h7a78: y = 16'h200;
			16'h7a79: y = 16'h200;
			16'h7a7a: y = 16'h200;
			16'h7a7b: y = 16'h200;
			16'h7a7c: y = 16'h200;
			16'h7a7d: y = 16'h200;
			16'h7a7e: y = 16'h200;
			16'h7a7f: y = 16'h200;
			16'h7a80: y = 16'h200;
			16'h7a81: y = 16'h200;
			16'h7a82: y = 16'h200;
			16'h7a83: y = 16'h200;
			16'h7a84: y = 16'h200;
			16'h7a85: y = 16'h200;
			16'h7a86: y = 16'h200;
			16'h7a87: y = 16'h200;
			16'h7a88: y = 16'h200;
			16'h7a89: y = 16'h200;
			16'h7a8a: y = 16'h200;
			16'h7a8b: y = 16'h200;
			16'h7a8c: y = 16'h200;
			16'h7a8d: y = 16'h200;
			16'h7a8e: y = 16'h200;
			16'h7a8f: y = 16'h200;
			16'h7a90: y = 16'h200;
			16'h7a91: y = 16'h200;
			16'h7a92: y = 16'h200;
			16'h7a93: y = 16'h200;
			16'h7a94: y = 16'h200;
			16'h7a95: y = 16'h200;
			16'h7a96: y = 16'h200;
			16'h7a97: y = 16'h200;
			16'h7a98: y = 16'h200;
			16'h7a99: y = 16'h200;
			16'h7a9a: y = 16'h200;
			16'h7a9b: y = 16'h200;
			16'h7a9c: y = 16'h200;
			16'h7a9d: y = 16'h200;
			16'h7a9e: y = 16'h200;
			16'h7a9f: y = 16'h200;
			16'h7aa0: y = 16'h200;
			16'h7aa1: y = 16'h200;
			16'h7aa2: y = 16'h200;
			16'h7aa3: y = 16'h200;
			16'h7aa4: y = 16'h200;
			16'h7aa5: y = 16'h200;
			16'h7aa6: y = 16'h200;
			16'h7aa7: y = 16'h200;
			16'h7aa8: y = 16'h200;
			16'h7aa9: y = 16'h200;
			16'h7aaa: y = 16'h200;
			16'h7aab: y = 16'h200;
			16'h7aac: y = 16'h200;
			16'h7aad: y = 16'h200;
			16'h7aae: y = 16'h200;
			16'h7aaf: y = 16'h200;
			16'h7ab0: y = 16'h200;
			16'h7ab1: y = 16'h200;
			16'h7ab2: y = 16'h200;
			16'h7ab3: y = 16'h200;
			16'h7ab4: y = 16'h200;
			16'h7ab5: y = 16'h200;
			16'h7ab6: y = 16'h200;
			16'h7ab7: y = 16'h200;
			16'h7ab8: y = 16'h200;
			16'h7ab9: y = 16'h200;
			16'h7aba: y = 16'h200;
			16'h7abb: y = 16'h200;
			16'h7abc: y = 16'h200;
			16'h7abd: y = 16'h200;
			16'h7abe: y = 16'h200;
			16'h7abf: y = 16'h200;
			16'h7ac0: y = 16'h200;
			16'h7ac1: y = 16'h200;
			16'h7ac2: y = 16'h200;
			16'h7ac3: y = 16'h200;
			16'h7ac4: y = 16'h200;
			16'h7ac5: y = 16'h200;
			16'h7ac6: y = 16'h200;
			16'h7ac7: y = 16'h200;
			16'h7ac8: y = 16'h200;
			16'h7ac9: y = 16'h200;
			16'h7aca: y = 16'h200;
			16'h7acb: y = 16'h200;
			16'h7acc: y = 16'h200;
			16'h7acd: y = 16'h200;
			16'h7ace: y = 16'h200;
			16'h7acf: y = 16'h200;
			16'h7ad0: y = 16'h200;
			16'h7ad1: y = 16'h200;
			16'h7ad2: y = 16'h200;
			16'h7ad3: y = 16'h200;
			16'h7ad4: y = 16'h200;
			16'h7ad5: y = 16'h200;
			16'h7ad6: y = 16'h200;
			16'h7ad7: y = 16'h200;
			16'h7ad8: y = 16'h200;
			16'h7ad9: y = 16'h200;
			16'h7ada: y = 16'h200;
			16'h7adb: y = 16'h200;
			16'h7adc: y = 16'h200;
			16'h7add: y = 16'h200;
			16'h7ade: y = 16'h200;
			16'h7adf: y = 16'h200;
			16'h7ae0: y = 16'h200;
			16'h7ae1: y = 16'h200;
			16'h7ae2: y = 16'h200;
			16'h7ae3: y = 16'h200;
			16'h7ae4: y = 16'h200;
			16'h7ae5: y = 16'h200;
			16'h7ae6: y = 16'h200;
			16'h7ae7: y = 16'h200;
			16'h7ae8: y = 16'h200;
			16'h7ae9: y = 16'h200;
			16'h7aea: y = 16'h200;
			16'h7aeb: y = 16'h200;
			16'h7aec: y = 16'h200;
			16'h7aed: y = 16'h200;
			16'h7aee: y = 16'h200;
			16'h7aef: y = 16'h200;
			16'h7af0: y = 16'h200;
			16'h7af1: y = 16'h200;
			16'h7af2: y = 16'h200;
			16'h7af3: y = 16'h200;
			16'h7af4: y = 16'h200;
			16'h7af5: y = 16'h200;
			16'h7af6: y = 16'h200;
			16'h7af7: y = 16'h200;
			16'h7af8: y = 16'h200;
			16'h7af9: y = 16'h200;
			16'h7afa: y = 16'h200;
			16'h7afb: y = 16'h200;
			16'h7afc: y = 16'h200;
			16'h7afd: y = 16'h200;
			16'h7afe: y = 16'h200;
			16'h7aff: y = 16'h200;
			16'h7b00: y = 16'h200;
			16'h7b01: y = 16'h200;
			16'h7b02: y = 16'h200;
			16'h7b03: y = 16'h200;
			16'h7b04: y = 16'h200;
			16'h7b05: y = 16'h200;
			16'h7b06: y = 16'h200;
			16'h7b07: y = 16'h200;
			16'h7b08: y = 16'h200;
			16'h7b09: y = 16'h200;
			16'h7b0a: y = 16'h200;
			16'h7b0b: y = 16'h200;
			16'h7b0c: y = 16'h200;
			16'h7b0d: y = 16'h200;
			16'h7b0e: y = 16'h200;
			16'h7b0f: y = 16'h200;
			16'h7b10: y = 16'h200;
			16'h7b11: y = 16'h200;
			16'h7b12: y = 16'h200;
			16'h7b13: y = 16'h200;
			16'h7b14: y = 16'h200;
			16'h7b15: y = 16'h200;
			16'h7b16: y = 16'h200;
			16'h7b17: y = 16'h200;
			16'h7b18: y = 16'h200;
			16'h7b19: y = 16'h200;
			16'h7b1a: y = 16'h200;
			16'h7b1b: y = 16'h200;
			16'h7b1c: y = 16'h200;
			16'h7b1d: y = 16'h200;
			16'h7b1e: y = 16'h200;
			16'h7b1f: y = 16'h200;
			16'h7b20: y = 16'h200;
			16'h7b21: y = 16'h200;
			16'h7b22: y = 16'h200;
			16'h7b23: y = 16'h200;
			16'h7b24: y = 16'h200;
			16'h7b25: y = 16'h200;
			16'h7b26: y = 16'h200;
			16'h7b27: y = 16'h200;
			16'h7b28: y = 16'h200;
			16'h7b29: y = 16'h200;
			16'h7b2a: y = 16'h200;
			16'h7b2b: y = 16'h200;
			16'h7b2c: y = 16'h200;
			16'h7b2d: y = 16'h200;
			16'h7b2e: y = 16'h200;
			16'h7b2f: y = 16'h200;
			16'h7b30: y = 16'h200;
			16'h7b31: y = 16'h200;
			16'h7b32: y = 16'h200;
			16'h7b33: y = 16'h200;
			16'h7b34: y = 16'h200;
			16'h7b35: y = 16'h200;
			16'h7b36: y = 16'h200;
			16'h7b37: y = 16'h200;
			16'h7b38: y = 16'h200;
			16'h7b39: y = 16'h200;
			16'h7b3a: y = 16'h200;
			16'h7b3b: y = 16'h200;
			16'h7b3c: y = 16'h200;
			16'h7b3d: y = 16'h200;
			16'h7b3e: y = 16'h200;
			16'h7b3f: y = 16'h200;
			16'h7b40: y = 16'h200;
			16'h7b41: y = 16'h200;
			16'h7b42: y = 16'h200;
			16'h7b43: y = 16'h200;
			16'h7b44: y = 16'h200;
			16'h7b45: y = 16'h200;
			16'h7b46: y = 16'h200;
			16'h7b47: y = 16'h200;
			16'h7b48: y = 16'h200;
			16'h7b49: y = 16'h200;
			16'h7b4a: y = 16'h200;
			16'h7b4b: y = 16'h200;
			16'h7b4c: y = 16'h200;
			16'h7b4d: y = 16'h200;
			16'h7b4e: y = 16'h200;
			16'h7b4f: y = 16'h200;
			16'h7b50: y = 16'h200;
			16'h7b51: y = 16'h200;
			16'h7b52: y = 16'h200;
			16'h7b53: y = 16'h200;
			16'h7b54: y = 16'h200;
			16'h7b55: y = 16'h200;
			16'h7b56: y = 16'h200;
			16'h7b57: y = 16'h200;
			16'h7b58: y = 16'h200;
			16'h7b59: y = 16'h200;
			16'h7b5a: y = 16'h200;
			16'h7b5b: y = 16'h200;
			16'h7b5c: y = 16'h200;
			16'h7b5d: y = 16'h200;
			16'h7b5e: y = 16'h200;
			16'h7b5f: y = 16'h200;
			16'h7b60: y = 16'h200;
			16'h7b61: y = 16'h200;
			16'h7b62: y = 16'h200;
			16'h7b63: y = 16'h200;
			16'h7b64: y = 16'h200;
			16'h7b65: y = 16'h200;
			16'h7b66: y = 16'h200;
			16'h7b67: y = 16'h200;
			16'h7b68: y = 16'h200;
			16'h7b69: y = 16'h200;
			16'h7b6a: y = 16'h200;
			16'h7b6b: y = 16'h200;
			16'h7b6c: y = 16'h200;
			16'h7b6d: y = 16'h200;
			16'h7b6e: y = 16'h200;
			16'h7b6f: y = 16'h200;
			16'h7b70: y = 16'h200;
			16'h7b71: y = 16'h200;
			16'h7b72: y = 16'h200;
			16'h7b73: y = 16'h200;
			16'h7b74: y = 16'h200;
			16'h7b75: y = 16'h200;
			16'h7b76: y = 16'h200;
			16'h7b77: y = 16'h200;
			16'h7b78: y = 16'h200;
			16'h7b79: y = 16'h200;
			16'h7b7a: y = 16'h200;
			16'h7b7b: y = 16'h200;
			16'h7b7c: y = 16'h200;
			16'h7b7d: y = 16'h200;
			16'h7b7e: y = 16'h200;
			16'h7b7f: y = 16'h200;
			16'h7b80: y = 16'h200;
			16'h7b81: y = 16'h200;
			16'h7b82: y = 16'h200;
			16'h7b83: y = 16'h200;
			16'h7b84: y = 16'h200;
			16'h7b85: y = 16'h200;
			16'h7b86: y = 16'h200;
			16'h7b87: y = 16'h200;
			16'h7b88: y = 16'h200;
			16'h7b89: y = 16'h200;
			16'h7b8a: y = 16'h200;
			16'h7b8b: y = 16'h200;
			16'h7b8c: y = 16'h200;
			16'h7b8d: y = 16'h200;
			16'h7b8e: y = 16'h200;
			16'h7b8f: y = 16'h200;
			16'h7b90: y = 16'h200;
			16'h7b91: y = 16'h200;
			16'h7b92: y = 16'h200;
			16'h7b93: y = 16'h200;
			16'h7b94: y = 16'h200;
			16'h7b95: y = 16'h200;
			16'h7b96: y = 16'h200;
			16'h7b97: y = 16'h200;
			16'h7b98: y = 16'h200;
			16'h7b99: y = 16'h200;
			16'h7b9a: y = 16'h200;
			16'h7b9b: y = 16'h200;
			16'h7b9c: y = 16'h200;
			16'h7b9d: y = 16'h200;
			16'h7b9e: y = 16'h200;
			16'h7b9f: y = 16'h200;
			16'h7ba0: y = 16'h200;
			16'h7ba1: y = 16'h200;
			16'h7ba2: y = 16'h200;
			16'h7ba3: y = 16'h200;
			16'h7ba4: y = 16'h200;
			16'h7ba5: y = 16'h200;
			16'h7ba6: y = 16'h200;
			16'h7ba7: y = 16'h200;
			16'h7ba8: y = 16'h200;
			16'h7ba9: y = 16'h200;
			16'h7baa: y = 16'h200;
			16'h7bab: y = 16'h200;
			16'h7bac: y = 16'h200;
			16'h7bad: y = 16'h200;
			16'h7bae: y = 16'h200;
			16'h7baf: y = 16'h200;
			16'h7bb0: y = 16'h200;
			16'h7bb1: y = 16'h200;
			16'h7bb2: y = 16'h200;
			16'h7bb3: y = 16'h200;
			16'h7bb4: y = 16'h200;
			16'h7bb5: y = 16'h200;
			16'h7bb6: y = 16'h200;
			16'h7bb7: y = 16'h200;
			16'h7bb8: y = 16'h200;
			16'h7bb9: y = 16'h200;
			16'h7bba: y = 16'h200;
			16'h7bbb: y = 16'h200;
			16'h7bbc: y = 16'h200;
			16'h7bbd: y = 16'h200;
			16'h7bbe: y = 16'h200;
			16'h7bbf: y = 16'h200;
			16'h7bc0: y = 16'h200;
			16'h7bc1: y = 16'h200;
			16'h7bc2: y = 16'h200;
			16'h7bc3: y = 16'h200;
			16'h7bc4: y = 16'h200;
			16'h7bc5: y = 16'h200;
			16'h7bc6: y = 16'h200;
			16'h7bc7: y = 16'h200;
			16'h7bc8: y = 16'h200;
			16'h7bc9: y = 16'h200;
			16'h7bca: y = 16'h200;
			16'h7bcb: y = 16'h200;
			16'h7bcc: y = 16'h200;
			16'h7bcd: y = 16'h200;
			16'h7bce: y = 16'h200;
			16'h7bcf: y = 16'h200;
			16'h7bd0: y = 16'h200;
			16'h7bd1: y = 16'h200;
			16'h7bd2: y = 16'h200;
			16'h7bd3: y = 16'h200;
			16'h7bd4: y = 16'h200;
			16'h7bd5: y = 16'h200;
			16'h7bd6: y = 16'h200;
			16'h7bd7: y = 16'h200;
			16'h7bd8: y = 16'h200;
			16'h7bd9: y = 16'h200;
			16'h7bda: y = 16'h200;
			16'h7bdb: y = 16'h200;
			16'h7bdc: y = 16'h200;
			16'h7bdd: y = 16'h200;
			16'h7bde: y = 16'h200;
			16'h7bdf: y = 16'h200;
			16'h7be0: y = 16'h200;
			16'h7be1: y = 16'h200;
			16'h7be2: y = 16'h200;
			16'h7be3: y = 16'h200;
			16'h7be4: y = 16'h200;
			16'h7be5: y = 16'h200;
			16'h7be6: y = 16'h200;
			16'h7be7: y = 16'h200;
			16'h7be8: y = 16'h200;
			16'h7be9: y = 16'h200;
			16'h7bea: y = 16'h200;
			16'h7beb: y = 16'h200;
			16'h7bec: y = 16'h200;
			16'h7bed: y = 16'h200;
			16'h7bee: y = 16'h200;
			16'h7bef: y = 16'h200;
			16'h7bf0: y = 16'h200;
			16'h7bf1: y = 16'h200;
			16'h7bf2: y = 16'h200;
			16'h7bf3: y = 16'h200;
			16'h7bf4: y = 16'h200;
			16'h7bf5: y = 16'h200;
			16'h7bf6: y = 16'h200;
			16'h7bf7: y = 16'h200;
			16'h7bf8: y = 16'h200;
			16'h7bf9: y = 16'h200;
			16'h7bfa: y = 16'h200;
			16'h7bfb: y = 16'h200;
			16'h7bfc: y = 16'h200;
			16'h7bfd: y = 16'h200;
			16'h7bfe: y = 16'h200;
			16'h7bff: y = 16'h200;
			16'h7c00: y = 16'h200;
			16'h7c01: y = 16'h200;
			16'h7c02: y = 16'h200;
			16'h7c03: y = 16'h200;
			16'h7c04: y = 16'h200;
			16'h7c05: y = 16'h200;
			16'h7c06: y = 16'h200;
			16'h7c07: y = 16'h200;
			16'h7c08: y = 16'h200;
			16'h7c09: y = 16'h200;
			16'h7c0a: y = 16'h200;
			16'h7c0b: y = 16'h200;
			16'h7c0c: y = 16'h200;
			16'h7c0d: y = 16'h200;
			16'h7c0e: y = 16'h200;
			16'h7c0f: y = 16'h200;
			16'h7c10: y = 16'h200;
			16'h7c11: y = 16'h200;
			16'h7c12: y = 16'h200;
			16'h7c13: y = 16'h200;
			16'h7c14: y = 16'h200;
			16'h7c15: y = 16'h200;
			16'h7c16: y = 16'h200;
			16'h7c17: y = 16'h200;
			16'h7c18: y = 16'h200;
			16'h7c19: y = 16'h200;
			16'h7c1a: y = 16'h200;
			16'h7c1b: y = 16'h200;
			16'h7c1c: y = 16'h200;
			16'h7c1d: y = 16'h200;
			16'h7c1e: y = 16'h200;
			16'h7c1f: y = 16'h200;
			16'h7c20: y = 16'h200;
			16'h7c21: y = 16'h200;
			16'h7c22: y = 16'h200;
			16'h7c23: y = 16'h200;
			16'h7c24: y = 16'h200;
			16'h7c25: y = 16'h200;
			16'h7c26: y = 16'h200;
			16'h7c27: y = 16'h200;
			16'h7c28: y = 16'h200;
			16'h7c29: y = 16'h200;
			16'h7c2a: y = 16'h200;
			16'h7c2b: y = 16'h200;
			16'h7c2c: y = 16'h200;
			16'h7c2d: y = 16'h200;
			16'h7c2e: y = 16'h200;
			16'h7c2f: y = 16'h200;
			16'h7c30: y = 16'h200;
			16'h7c31: y = 16'h200;
			16'h7c32: y = 16'h200;
			16'h7c33: y = 16'h200;
			16'h7c34: y = 16'h200;
			16'h7c35: y = 16'h200;
			16'h7c36: y = 16'h200;
			16'h7c37: y = 16'h200;
			16'h7c38: y = 16'h200;
			16'h7c39: y = 16'h200;
			16'h7c3a: y = 16'h200;
			16'h7c3b: y = 16'h200;
			16'h7c3c: y = 16'h200;
			16'h7c3d: y = 16'h200;
			16'h7c3e: y = 16'h200;
			16'h7c3f: y = 16'h200;
			16'h7c40: y = 16'h200;
			16'h7c41: y = 16'h200;
			16'h7c42: y = 16'h200;
			16'h7c43: y = 16'h200;
			16'h7c44: y = 16'h200;
			16'h7c45: y = 16'h200;
			16'h7c46: y = 16'h200;
			16'h7c47: y = 16'h200;
			16'h7c48: y = 16'h200;
			16'h7c49: y = 16'h200;
			16'h7c4a: y = 16'h200;
			16'h7c4b: y = 16'h200;
			16'h7c4c: y = 16'h200;
			16'h7c4d: y = 16'h200;
			16'h7c4e: y = 16'h200;
			16'h7c4f: y = 16'h200;
			16'h7c50: y = 16'h200;
			16'h7c51: y = 16'h200;
			16'h7c52: y = 16'h200;
			16'h7c53: y = 16'h200;
			16'h7c54: y = 16'h200;
			16'h7c55: y = 16'h200;
			16'h7c56: y = 16'h200;
			16'h7c57: y = 16'h200;
			16'h7c58: y = 16'h200;
			16'h7c59: y = 16'h200;
			16'h7c5a: y = 16'h200;
			16'h7c5b: y = 16'h200;
			16'h7c5c: y = 16'h200;
			16'h7c5d: y = 16'h200;
			16'h7c5e: y = 16'h200;
			16'h7c5f: y = 16'h200;
			16'h7c60: y = 16'h200;
			16'h7c61: y = 16'h200;
			16'h7c62: y = 16'h200;
			16'h7c63: y = 16'h200;
			16'h7c64: y = 16'h200;
			16'h7c65: y = 16'h200;
			16'h7c66: y = 16'h200;
			16'h7c67: y = 16'h200;
			16'h7c68: y = 16'h200;
			16'h7c69: y = 16'h200;
			16'h7c6a: y = 16'h200;
			16'h7c6b: y = 16'h200;
			16'h7c6c: y = 16'h200;
			16'h7c6d: y = 16'h200;
			16'h7c6e: y = 16'h200;
			16'h7c6f: y = 16'h200;
			16'h7c70: y = 16'h200;
			16'h7c71: y = 16'h200;
			16'h7c72: y = 16'h200;
			16'h7c73: y = 16'h200;
			16'h7c74: y = 16'h200;
			16'h7c75: y = 16'h200;
			16'h7c76: y = 16'h200;
			16'h7c77: y = 16'h200;
			16'h7c78: y = 16'h200;
			16'h7c79: y = 16'h200;
			16'h7c7a: y = 16'h200;
			16'h7c7b: y = 16'h200;
			16'h7c7c: y = 16'h200;
			16'h7c7d: y = 16'h200;
			16'h7c7e: y = 16'h200;
			16'h7c7f: y = 16'h200;
			16'h7c80: y = 16'h200;
			16'h7c81: y = 16'h200;
			16'h7c82: y = 16'h200;
			16'h7c83: y = 16'h200;
			16'h7c84: y = 16'h200;
			16'h7c85: y = 16'h200;
			16'h7c86: y = 16'h200;
			16'h7c87: y = 16'h200;
			16'h7c88: y = 16'h200;
			16'h7c89: y = 16'h200;
			16'h7c8a: y = 16'h200;
			16'h7c8b: y = 16'h200;
			16'h7c8c: y = 16'h200;
			16'h7c8d: y = 16'h200;
			16'h7c8e: y = 16'h200;
			16'h7c8f: y = 16'h200;
			16'h7c90: y = 16'h200;
			16'h7c91: y = 16'h200;
			16'h7c92: y = 16'h200;
			16'h7c93: y = 16'h200;
			16'h7c94: y = 16'h200;
			16'h7c95: y = 16'h200;
			16'h7c96: y = 16'h200;
			16'h7c97: y = 16'h200;
			16'h7c98: y = 16'h200;
			16'h7c99: y = 16'h200;
			16'h7c9a: y = 16'h200;
			16'h7c9b: y = 16'h200;
			16'h7c9c: y = 16'h200;
			16'h7c9d: y = 16'h200;
			16'h7c9e: y = 16'h200;
			16'h7c9f: y = 16'h200;
			16'h7ca0: y = 16'h200;
			16'h7ca1: y = 16'h200;
			16'h7ca2: y = 16'h200;
			16'h7ca3: y = 16'h200;
			16'h7ca4: y = 16'h200;
			16'h7ca5: y = 16'h200;
			16'h7ca6: y = 16'h200;
			16'h7ca7: y = 16'h200;
			16'h7ca8: y = 16'h200;
			16'h7ca9: y = 16'h200;
			16'h7caa: y = 16'h200;
			16'h7cab: y = 16'h200;
			16'h7cac: y = 16'h200;
			16'h7cad: y = 16'h200;
			16'h7cae: y = 16'h200;
			16'h7caf: y = 16'h200;
			16'h7cb0: y = 16'h200;
			16'h7cb1: y = 16'h200;
			16'h7cb2: y = 16'h200;
			16'h7cb3: y = 16'h200;
			16'h7cb4: y = 16'h200;
			16'h7cb5: y = 16'h200;
			16'h7cb6: y = 16'h200;
			16'h7cb7: y = 16'h200;
			16'h7cb8: y = 16'h200;
			16'h7cb9: y = 16'h200;
			16'h7cba: y = 16'h200;
			16'h7cbb: y = 16'h200;
			16'h7cbc: y = 16'h200;
			16'h7cbd: y = 16'h200;
			16'h7cbe: y = 16'h200;
			16'h7cbf: y = 16'h200;
			16'h7cc0: y = 16'h200;
			16'h7cc1: y = 16'h200;
			16'h7cc2: y = 16'h200;
			16'h7cc3: y = 16'h200;
			16'h7cc4: y = 16'h200;
			16'h7cc5: y = 16'h200;
			16'h7cc6: y = 16'h200;
			16'h7cc7: y = 16'h200;
			16'h7cc8: y = 16'h200;
			16'h7cc9: y = 16'h200;
			16'h7cca: y = 16'h200;
			16'h7ccb: y = 16'h200;
			16'h7ccc: y = 16'h200;
			16'h7ccd: y = 16'h200;
			16'h7cce: y = 16'h200;
			16'h7ccf: y = 16'h200;
			16'h7cd0: y = 16'h200;
			16'h7cd1: y = 16'h200;
			16'h7cd2: y = 16'h200;
			16'h7cd3: y = 16'h200;
			16'h7cd4: y = 16'h200;
			16'h7cd5: y = 16'h200;
			16'h7cd6: y = 16'h200;
			16'h7cd7: y = 16'h200;
			16'h7cd8: y = 16'h200;
			16'h7cd9: y = 16'h200;
			16'h7cda: y = 16'h200;
			16'h7cdb: y = 16'h200;
			16'h7cdc: y = 16'h200;
			16'h7cdd: y = 16'h200;
			16'h7cde: y = 16'h200;
			16'h7cdf: y = 16'h200;
			16'h7ce0: y = 16'h200;
			16'h7ce1: y = 16'h200;
			16'h7ce2: y = 16'h200;
			16'h7ce3: y = 16'h200;
			16'h7ce4: y = 16'h200;
			16'h7ce5: y = 16'h200;
			16'h7ce6: y = 16'h200;
			16'h7ce7: y = 16'h200;
			16'h7ce8: y = 16'h200;
			16'h7ce9: y = 16'h200;
			16'h7cea: y = 16'h200;
			16'h7ceb: y = 16'h200;
			16'h7cec: y = 16'h200;
			16'h7ced: y = 16'h200;
			16'h7cee: y = 16'h200;
			16'h7cef: y = 16'h200;
			16'h7cf0: y = 16'h200;
			16'h7cf1: y = 16'h200;
			16'h7cf2: y = 16'h200;
			16'h7cf3: y = 16'h200;
			16'h7cf4: y = 16'h200;
			16'h7cf5: y = 16'h200;
			16'h7cf6: y = 16'h200;
			16'h7cf7: y = 16'h200;
			16'h7cf8: y = 16'h200;
			16'h7cf9: y = 16'h200;
			16'h7cfa: y = 16'h200;
			16'h7cfb: y = 16'h200;
			16'h7cfc: y = 16'h200;
			16'h7cfd: y = 16'h200;
			16'h7cfe: y = 16'h200;
			16'h7cff: y = 16'h200;
			16'h7d00: y = 16'h200;
			16'h7d01: y = 16'h200;
			16'h7d02: y = 16'h200;
			16'h7d03: y = 16'h200;
			16'h7d04: y = 16'h200;
			16'h7d05: y = 16'h200;
			16'h7d06: y = 16'h200;
			16'h7d07: y = 16'h200;
			16'h7d08: y = 16'h200;
			16'h7d09: y = 16'h200;
			16'h7d0a: y = 16'h200;
			16'h7d0b: y = 16'h200;
			16'h7d0c: y = 16'h200;
			16'h7d0d: y = 16'h200;
			16'h7d0e: y = 16'h200;
			16'h7d0f: y = 16'h200;
			16'h7d10: y = 16'h200;
			16'h7d11: y = 16'h200;
			16'h7d12: y = 16'h200;
			16'h7d13: y = 16'h200;
			16'h7d14: y = 16'h200;
			16'h7d15: y = 16'h200;
			16'h7d16: y = 16'h200;
			16'h7d17: y = 16'h200;
			16'h7d18: y = 16'h200;
			16'h7d19: y = 16'h200;
			16'h7d1a: y = 16'h200;
			16'h7d1b: y = 16'h200;
			16'h7d1c: y = 16'h200;
			16'h7d1d: y = 16'h200;
			16'h7d1e: y = 16'h200;
			16'h7d1f: y = 16'h200;
			16'h7d20: y = 16'h200;
			16'h7d21: y = 16'h200;
			16'h7d22: y = 16'h200;
			16'h7d23: y = 16'h200;
			16'h7d24: y = 16'h200;
			16'h7d25: y = 16'h200;
			16'h7d26: y = 16'h200;
			16'h7d27: y = 16'h200;
			16'h7d28: y = 16'h200;
			16'h7d29: y = 16'h200;
			16'h7d2a: y = 16'h200;
			16'h7d2b: y = 16'h200;
			16'h7d2c: y = 16'h200;
			16'h7d2d: y = 16'h200;
			16'h7d2e: y = 16'h200;
			16'h7d2f: y = 16'h200;
			16'h7d30: y = 16'h200;
			16'h7d31: y = 16'h200;
			16'h7d32: y = 16'h200;
			16'h7d33: y = 16'h200;
			16'h7d34: y = 16'h200;
			16'h7d35: y = 16'h200;
			16'h7d36: y = 16'h200;
			16'h7d37: y = 16'h200;
			16'h7d38: y = 16'h200;
			16'h7d39: y = 16'h200;
			16'h7d3a: y = 16'h200;
			16'h7d3b: y = 16'h200;
			16'h7d3c: y = 16'h200;
			16'h7d3d: y = 16'h200;
			16'h7d3e: y = 16'h200;
			16'h7d3f: y = 16'h200;
			16'h7d40: y = 16'h200;
			16'h7d41: y = 16'h200;
			16'h7d42: y = 16'h200;
			16'h7d43: y = 16'h200;
			16'h7d44: y = 16'h200;
			16'h7d45: y = 16'h200;
			16'h7d46: y = 16'h200;
			16'h7d47: y = 16'h200;
			16'h7d48: y = 16'h200;
			16'h7d49: y = 16'h200;
			16'h7d4a: y = 16'h200;
			16'h7d4b: y = 16'h200;
			16'h7d4c: y = 16'h200;
			16'h7d4d: y = 16'h200;
			16'h7d4e: y = 16'h200;
			16'h7d4f: y = 16'h200;
			16'h7d50: y = 16'h200;
			16'h7d51: y = 16'h200;
			16'h7d52: y = 16'h200;
			16'h7d53: y = 16'h200;
			16'h7d54: y = 16'h200;
			16'h7d55: y = 16'h200;
			16'h7d56: y = 16'h200;
			16'h7d57: y = 16'h200;
			16'h7d58: y = 16'h200;
			16'h7d59: y = 16'h200;
			16'h7d5a: y = 16'h200;
			16'h7d5b: y = 16'h200;
			16'h7d5c: y = 16'h200;
			16'h7d5d: y = 16'h200;
			16'h7d5e: y = 16'h200;
			16'h7d5f: y = 16'h200;
			16'h7d60: y = 16'h200;
			16'h7d61: y = 16'h200;
			16'h7d62: y = 16'h200;
			16'h7d63: y = 16'h200;
			16'h7d64: y = 16'h200;
			16'h7d65: y = 16'h200;
			16'h7d66: y = 16'h200;
			16'h7d67: y = 16'h200;
			16'h7d68: y = 16'h200;
			16'h7d69: y = 16'h200;
			16'h7d6a: y = 16'h200;
			16'h7d6b: y = 16'h200;
			16'h7d6c: y = 16'h200;
			16'h7d6d: y = 16'h200;
			16'h7d6e: y = 16'h200;
			16'h7d6f: y = 16'h200;
			16'h7d70: y = 16'h200;
			16'h7d71: y = 16'h200;
			16'h7d72: y = 16'h200;
			16'h7d73: y = 16'h200;
			16'h7d74: y = 16'h200;
			16'h7d75: y = 16'h200;
			16'h7d76: y = 16'h200;
			16'h7d77: y = 16'h200;
			16'h7d78: y = 16'h200;
			16'h7d79: y = 16'h200;
			16'h7d7a: y = 16'h200;
			16'h7d7b: y = 16'h200;
			16'h7d7c: y = 16'h200;
			16'h7d7d: y = 16'h200;
			16'h7d7e: y = 16'h200;
			16'h7d7f: y = 16'h200;
			16'h7d80: y = 16'h200;
			16'h7d81: y = 16'h200;
			16'h7d82: y = 16'h200;
			16'h7d83: y = 16'h200;
			16'h7d84: y = 16'h200;
			16'h7d85: y = 16'h200;
			16'h7d86: y = 16'h200;
			16'h7d87: y = 16'h200;
			16'h7d88: y = 16'h200;
			16'h7d89: y = 16'h200;
			16'h7d8a: y = 16'h200;
			16'h7d8b: y = 16'h200;
			16'h7d8c: y = 16'h200;
			16'h7d8d: y = 16'h200;
			16'h7d8e: y = 16'h200;
			16'h7d8f: y = 16'h200;
			16'h7d90: y = 16'h200;
			16'h7d91: y = 16'h200;
			16'h7d92: y = 16'h200;
			16'h7d93: y = 16'h200;
			16'h7d94: y = 16'h200;
			16'h7d95: y = 16'h200;
			16'h7d96: y = 16'h200;
			16'h7d97: y = 16'h200;
			16'h7d98: y = 16'h200;
			16'h7d99: y = 16'h200;
			16'h7d9a: y = 16'h200;
			16'h7d9b: y = 16'h200;
			16'h7d9c: y = 16'h200;
			16'h7d9d: y = 16'h200;
			16'h7d9e: y = 16'h200;
			16'h7d9f: y = 16'h200;
			16'h7da0: y = 16'h200;
			16'h7da1: y = 16'h200;
			16'h7da2: y = 16'h200;
			16'h7da3: y = 16'h200;
			16'h7da4: y = 16'h200;
			16'h7da5: y = 16'h200;
			16'h7da6: y = 16'h200;
			16'h7da7: y = 16'h200;
			16'h7da8: y = 16'h200;
			16'h7da9: y = 16'h200;
			16'h7daa: y = 16'h200;
			16'h7dab: y = 16'h200;
			16'h7dac: y = 16'h200;
			16'h7dad: y = 16'h200;
			16'h7dae: y = 16'h200;
			16'h7daf: y = 16'h200;
			16'h7db0: y = 16'h200;
			16'h7db1: y = 16'h200;
			16'h7db2: y = 16'h200;
			16'h7db3: y = 16'h200;
			16'h7db4: y = 16'h200;
			16'h7db5: y = 16'h200;
			16'h7db6: y = 16'h200;
			16'h7db7: y = 16'h200;
			16'h7db8: y = 16'h200;
			16'h7db9: y = 16'h200;
			16'h7dba: y = 16'h200;
			16'h7dbb: y = 16'h200;
			16'h7dbc: y = 16'h200;
			16'h7dbd: y = 16'h200;
			16'h7dbe: y = 16'h200;
			16'h7dbf: y = 16'h200;
			16'h7dc0: y = 16'h200;
			16'h7dc1: y = 16'h200;
			16'h7dc2: y = 16'h200;
			16'h7dc3: y = 16'h200;
			16'h7dc4: y = 16'h200;
			16'h7dc5: y = 16'h200;
			16'h7dc6: y = 16'h200;
			16'h7dc7: y = 16'h200;
			16'h7dc8: y = 16'h200;
			16'h7dc9: y = 16'h200;
			16'h7dca: y = 16'h200;
			16'h7dcb: y = 16'h200;
			16'h7dcc: y = 16'h200;
			16'h7dcd: y = 16'h200;
			16'h7dce: y = 16'h200;
			16'h7dcf: y = 16'h200;
			16'h7dd0: y = 16'h200;
			16'h7dd1: y = 16'h200;
			16'h7dd2: y = 16'h200;
			16'h7dd3: y = 16'h200;
			16'h7dd4: y = 16'h200;
			16'h7dd5: y = 16'h200;
			16'h7dd6: y = 16'h200;
			16'h7dd7: y = 16'h200;
			16'h7dd8: y = 16'h200;
			16'h7dd9: y = 16'h200;
			16'h7dda: y = 16'h200;
			16'h7ddb: y = 16'h200;
			16'h7ddc: y = 16'h200;
			16'h7ddd: y = 16'h200;
			16'h7dde: y = 16'h200;
			16'h7ddf: y = 16'h200;
			16'h7de0: y = 16'h200;
			16'h7de1: y = 16'h200;
			16'h7de2: y = 16'h200;
			16'h7de3: y = 16'h200;
			16'h7de4: y = 16'h200;
			16'h7de5: y = 16'h200;
			16'h7de6: y = 16'h200;
			16'h7de7: y = 16'h200;
			16'h7de8: y = 16'h200;
			16'h7de9: y = 16'h200;
			16'h7dea: y = 16'h200;
			16'h7deb: y = 16'h200;
			16'h7dec: y = 16'h200;
			16'h7ded: y = 16'h200;
			16'h7dee: y = 16'h200;
			16'h7def: y = 16'h200;
			16'h7df0: y = 16'h200;
			16'h7df1: y = 16'h200;
			16'h7df2: y = 16'h200;
			16'h7df3: y = 16'h200;
			16'h7df4: y = 16'h200;
			16'h7df5: y = 16'h200;
			16'h7df6: y = 16'h200;
			16'h7df7: y = 16'h200;
			16'h7df8: y = 16'h200;
			16'h7df9: y = 16'h200;
			16'h7dfa: y = 16'h200;
			16'h7dfb: y = 16'h200;
			16'h7dfc: y = 16'h200;
			16'h7dfd: y = 16'h200;
			16'h7dfe: y = 16'h200;
			16'h7dff: y = 16'h200;
			16'h7e00: y = 16'h200;
			16'h7e01: y = 16'h200;
			16'h7e02: y = 16'h200;
			16'h7e03: y = 16'h200;
			16'h7e04: y = 16'h200;
			16'h7e05: y = 16'h200;
			16'h7e06: y = 16'h200;
			16'h7e07: y = 16'h200;
			16'h7e08: y = 16'h200;
			16'h7e09: y = 16'h200;
			16'h7e0a: y = 16'h200;
			16'h7e0b: y = 16'h200;
			16'h7e0c: y = 16'h200;
			16'h7e0d: y = 16'h200;
			16'h7e0e: y = 16'h200;
			16'h7e0f: y = 16'h200;
			16'h7e10: y = 16'h200;
			16'h7e11: y = 16'h200;
			16'h7e12: y = 16'h200;
			16'h7e13: y = 16'h200;
			16'h7e14: y = 16'h200;
			16'h7e15: y = 16'h200;
			16'h7e16: y = 16'h200;
			16'h7e17: y = 16'h200;
			16'h7e18: y = 16'h200;
			16'h7e19: y = 16'h200;
			16'h7e1a: y = 16'h200;
			16'h7e1b: y = 16'h200;
			16'h7e1c: y = 16'h200;
			16'h7e1d: y = 16'h200;
			16'h7e1e: y = 16'h200;
			16'h7e1f: y = 16'h200;
			16'h7e20: y = 16'h200;
			16'h7e21: y = 16'h200;
			16'h7e22: y = 16'h200;
			16'h7e23: y = 16'h200;
			16'h7e24: y = 16'h200;
			16'h7e25: y = 16'h200;
			16'h7e26: y = 16'h200;
			16'h7e27: y = 16'h200;
			16'h7e28: y = 16'h200;
			16'h7e29: y = 16'h200;
			16'h7e2a: y = 16'h200;
			16'h7e2b: y = 16'h200;
			16'h7e2c: y = 16'h200;
			16'h7e2d: y = 16'h200;
			16'h7e2e: y = 16'h200;
			16'h7e2f: y = 16'h200;
			16'h7e30: y = 16'h200;
			16'h7e31: y = 16'h200;
			16'h7e32: y = 16'h200;
			16'h7e33: y = 16'h200;
			16'h7e34: y = 16'h200;
			16'h7e35: y = 16'h200;
			16'h7e36: y = 16'h200;
			16'h7e37: y = 16'h200;
			16'h7e38: y = 16'h200;
			16'h7e39: y = 16'h200;
			16'h7e3a: y = 16'h200;
			16'h7e3b: y = 16'h200;
			16'h7e3c: y = 16'h200;
			16'h7e3d: y = 16'h200;
			16'h7e3e: y = 16'h200;
			16'h7e3f: y = 16'h200;
			16'h7e40: y = 16'h200;
			16'h7e41: y = 16'h200;
			16'h7e42: y = 16'h200;
			16'h7e43: y = 16'h200;
			16'h7e44: y = 16'h200;
			16'h7e45: y = 16'h200;
			16'h7e46: y = 16'h200;
			16'h7e47: y = 16'h200;
			16'h7e48: y = 16'h200;
			16'h7e49: y = 16'h200;
			16'h7e4a: y = 16'h200;
			16'h7e4b: y = 16'h200;
			16'h7e4c: y = 16'h200;
			16'h7e4d: y = 16'h200;
			16'h7e4e: y = 16'h200;
			16'h7e4f: y = 16'h200;
			16'h7e50: y = 16'h200;
			16'h7e51: y = 16'h200;
			16'h7e52: y = 16'h200;
			16'h7e53: y = 16'h200;
			16'h7e54: y = 16'h200;
			16'h7e55: y = 16'h200;
			16'h7e56: y = 16'h200;
			16'h7e57: y = 16'h200;
			16'h7e58: y = 16'h200;
			16'h7e59: y = 16'h200;
			16'h7e5a: y = 16'h200;
			16'h7e5b: y = 16'h200;
			16'h7e5c: y = 16'h200;
			16'h7e5d: y = 16'h200;
			16'h7e5e: y = 16'h200;
			16'h7e5f: y = 16'h200;
			16'h7e60: y = 16'h200;
			16'h7e61: y = 16'h200;
			16'h7e62: y = 16'h200;
			16'h7e63: y = 16'h200;
			16'h7e64: y = 16'h200;
			16'h7e65: y = 16'h200;
			16'h7e66: y = 16'h200;
			16'h7e67: y = 16'h200;
			16'h7e68: y = 16'h200;
			16'h7e69: y = 16'h200;
			16'h7e6a: y = 16'h200;
			16'h7e6b: y = 16'h200;
			16'h7e6c: y = 16'h200;
			16'h7e6d: y = 16'h200;
			16'h7e6e: y = 16'h200;
			16'h7e6f: y = 16'h200;
			16'h7e70: y = 16'h200;
			16'h7e71: y = 16'h200;
			16'h7e72: y = 16'h200;
			16'h7e73: y = 16'h200;
			16'h7e74: y = 16'h200;
			16'h7e75: y = 16'h200;
			16'h7e76: y = 16'h200;
			16'h7e77: y = 16'h200;
			16'h7e78: y = 16'h200;
			16'h7e79: y = 16'h200;
			16'h7e7a: y = 16'h200;
			16'h7e7b: y = 16'h200;
			16'h7e7c: y = 16'h200;
			16'h7e7d: y = 16'h200;
			16'h7e7e: y = 16'h200;
			16'h7e7f: y = 16'h200;
			16'h7e80: y = 16'h200;
			16'h7e81: y = 16'h200;
			16'h7e82: y = 16'h200;
			16'h7e83: y = 16'h200;
			16'h7e84: y = 16'h200;
			16'h7e85: y = 16'h200;
			16'h7e86: y = 16'h200;
			16'h7e87: y = 16'h200;
			16'h7e88: y = 16'h200;
			16'h7e89: y = 16'h200;
			16'h7e8a: y = 16'h200;
			16'h7e8b: y = 16'h200;
			16'h7e8c: y = 16'h200;
			16'h7e8d: y = 16'h200;
			16'h7e8e: y = 16'h200;
			16'h7e8f: y = 16'h200;
			16'h7e90: y = 16'h200;
			16'h7e91: y = 16'h200;
			16'h7e92: y = 16'h200;
			16'h7e93: y = 16'h200;
			16'h7e94: y = 16'h200;
			16'h7e95: y = 16'h200;
			16'h7e96: y = 16'h200;
			16'h7e97: y = 16'h200;
			16'h7e98: y = 16'h200;
			16'h7e99: y = 16'h200;
			16'h7e9a: y = 16'h200;
			16'h7e9b: y = 16'h200;
			16'h7e9c: y = 16'h200;
			16'h7e9d: y = 16'h200;
			16'h7e9e: y = 16'h200;
			16'h7e9f: y = 16'h200;
			16'h7ea0: y = 16'h200;
			16'h7ea1: y = 16'h200;
			16'h7ea2: y = 16'h200;
			16'h7ea3: y = 16'h200;
			16'h7ea4: y = 16'h200;
			16'h7ea5: y = 16'h200;
			16'h7ea6: y = 16'h200;
			16'h7ea7: y = 16'h200;
			16'h7ea8: y = 16'h200;
			16'h7ea9: y = 16'h200;
			16'h7eaa: y = 16'h200;
			16'h7eab: y = 16'h200;
			16'h7eac: y = 16'h200;
			16'h7ead: y = 16'h200;
			16'h7eae: y = 16'h200;
			16'h7eaf: y = 16'h200;
			16'h7eb0: y = 16'h200;
			16'h7eb1: y = 16'h200;
			16'h7eb2: y = 16'h200;
			16'h7eb3: y = 16'h200;
			16'h7eb4: y = 16'h200;
			16'h7eb5: y = 16'h200;
			16'h7eb6: y = 16'h200;
			16'h7eb7: y = 16'h200;
			16'h7eb8: y = 16'h200;
			16'h7eb9: y = 16'h200;
			16'h7eba: y = 16'h200;
			16'h7ebb: y = 16'h200;
			16'h7ebc: y = 16'h200;
			16'h7ebd: y = 16'h200;
			16'h7ebe: y = 16'h200;
			16'h7ebf: y = 16'h200;
			16'h7ec0: y = 16'h200;
			16'h7ec1: y = 16'h200;
			16'h7ec2: y = 16'h200;
			16'h7ec3: y = 16'h200;
			16'h7ec4: y = 16'h200;
			16'h7ec5: y = 16'h200;
			16'h7ec6: y = 16'h200;
			16'h7ec7: y = 16'h200;
			16'h7ec8: y = 16'h200;
			16'h7ec9: y = 16'h200;
			16'h7eca: y = 16'h200;
			16'h7ecb: y = 16'h200;
			16'h7ecc: y = 16'h200;
			16'h7ecd: y = 16'h200;
			16'h7ece: y = 16'h200;
			16'h7ecf: y = 16'h200;
			16'h7ed0: y = 16'h200;
			16'h7ed1: y = 16'h200;
			16'h7ed2: y = 16'h200;
			16'h7ed3: y = 16'h200;
			16'h7ed4: y = 16'h200;
			16'h7ed5: y = 16'h200;
			16'h7ed6: y = 16'h200;
			16'h7ed7: y = 16'h200;
			16'h7ed8: y = 16'h200;
			16'h7ed9: y = 16'h200;
			16'h7eda: y = 16'h200;
			16'h7edb: y = 16'h200;
			16'h7edc: y = 16'h200;
			16'h7edd: y = 16'h200;
			16'h7ede: y = 16'h200;
			16'h7edf: y = 16'h200;
			16'h7ee0: y = 16'h200;
			16'h7ee1: y = 16'h200;
			16'h7ee2: y = 16'h200;
			16'h7ee3: y = 16'h200;
			16'h7ee4: y = 16'h200;
			16'h7ee5: y = 16'h200;
			16'h7ee6: y = 16'h200;
			16'h7ee7: y = 16'h200;
			16'h7ee8: y = 16'h200;
			16'h7ee9: y = 16'h200;
			16'h7eea: y = 16'h200;
			16'h7eeb: y = 16'h200;
			16'h7eec: y = 16'h200;
			16'h7eed: y = 16'h200;
			16'h7eee: y = 16'h200;
			16'h7eef: y = 16'h200;
			16'h7ef0: y = 16'h200;
			16'h7ef1: y = 16'h200;
			16'h7ef2: y = 16'h200;
			16'h7ef3: y = 16'h200;
			16'h7ef4: y = 16'h200;
			16'h7ef5: y = 16'h200;
			16'h7ef6: y = 16'h200;
			16'h7ef7: y = 16'h200;
			16'h7ef8: y = 16'h200;
			16'h7ef9: y = 16'h200;
			16'h7efa: y = 16'h200;
			16'h7efb: y = 16'h200;
			16'h7efc: y = 16'h200;
			16'h7efd: y = 16'h200;
			16'h7efe: y = 16'h200;
			16'h7eff: y = 16'h200;
			16'h7f00: y = 16'h200;
			16'h7f01: y = 16'h200;
			16'h7f02: y = 16'h200;
			16'h7f03: y = 16'h200;
			16'h7f04: y = 16'h200;
			16'h7f05: y = 16'h200;
			16'h7f06: y = 16'h200;
			16'h7f07: y = 16'h200;
			16'h7f08: y = 16'h200;
			16'h7f09: y = 16'h200;
			16'h7f0a: y = 16'h200;
			16'h7f0b: y = 16'h200;
			16'h7f0c: y = 16'h200;
			16'h7f0d: y = 16'h200;
			16'h7f0e: y = 16'h200;
			16'h7f0f: y = 16'h200;
			16'h7f10: y = 16'h200;
			16'h7f11: y = 16'h200;
			16'h7f12: y = 16'h200;
			16'h7f13: y = 16'h200;
			16'h7f14: y = 16'h200;
			16'h7f15: y = 16'h200;
			16'h7f16: y = 16'h200;
			16'h7f17: y = 16'h200;
			16'h7f18: y = 16'h200;
			16'h7f19: y = 16'h200;
			16'h7f1a: y = 16'h200;
			16'h7f1b: y = 16'h200;
			16'h7f1c: y = 16'h200;
			16'h7f1d: y = 16'h200;
			16'h7f1e: y = 16'h200;
			16'h7f1f: y = 16'h200;
			16'h7f20: y = 16'h200;
			16'h7f21: y = 16'h200;
			16'h7f22: y = 16'h200;
			16'h7f23: y = 16'h200;
			16'h7f24: y = 16'h200;
			16'h7f25: y = 16'h200;
			16'h7f26: y = 16'h200;
			16'h7f27: y = 16'h200;
			16'h7f28: y = 16'h200;
			16'h7f29: y = 16'h200;
			16'h7f2a: y = 16'h200;
			16'h7f2b: y = 16'h200;
			16'h7f2c: y = 16'h200;
			16'h7f2d: y = 16'h200;
			16'h7f2e: y = 16'h200;
			16'h7f2f: y = 16'h200;
			16'h7f30: y = 16'h200;
			16'h7f31: y = 16'h200;
			16'h7f32: y = 16'h200;
			16'h7f33: y = 16'h200;
			16'h7f34: y = 16'h200;
			16'h7f35: y = 16'h200;
			16'h7f36: y = 16'h200;
			16'h7f37: y = 16'h200;
			16'h7f38: y = 16'h200;
			16'h7f39: y = 16'h200;
			16'h7f3a: y = 16'h200;
			16'h7f3b: y = 16'h200;
			16'h7f3c: y = 16'h200;
			16'h7f3d: y = 16'h200;
			16'h7f3e: y = 16'h200;
			16'h7f3f: y = 16'h200;
			16'h7f40: y = 16'h200;
			16'h7f41: y = 16'h200;
			16'h7f42: y = 16'h200;
			16'h7f43: y = 16'h200;
			16'h7f44: y = 16'h200;
			16'h7f45: y = 16'h200;
			16'h7f46: y = 16'h200;
			16'h7f47: y = 16'h200;
			16'h7f48: y = 16'h200;
			16'h7f49: y = 16'h200;
			16'h7f4a: y = 16'h200;
			16'h7f4b: y = 16'h200;
			16'h7f4c: y = 16'h200;
			16'h7f4d: y = 16'h200;
			16'h7f4e: y = 16'h200;
			16'h7f4f: y = 16'h200;
			16'h7f50: y = 16'h200;
			16'h7f51: y = 16'h200;
			16'h7f52: y = 16'h200;
			16'h7f53: y = 16'h200;
			16'h7f54: y = 16'h200;
			16'h7f55: y = 16'h200;
			16'h7f56: y = 16'h200;
			16'h7f57: y = 16'h200;
			16'h7f58: y = 16'h200;
			16'h7f59: y = 16'h200;
			16'h7f5a: y = 16'h200;
			16'h7f5b: y = 16'h200;
			16'h7f5c: y = 16'h200;
			16'h7f5d: y = 16'h200;
			16'h7f5e: y = 16'h200;
			16'h7f5f: y = 16'h200;
			16'h7f60: y = 16'h200;
			16'h7f61: y = 16'h200;
			16'h7f62: y = 16'h200;
			16'h7f63: y = 16'h200;
			16'h7f64: y = 16'h200;
			16'h7f65: y = 16'h200;
			16'h7f66: y = 16'h200;
			16'h7f67: y = 16'h200;
			16'h7f68: y = 16'h200;
			16'h7f69: y = 16'h200;
			16'h7f6a: y = 16'h200;
			16'h7f6b: y = 16'h200;
			16'h7f6c: y = 16'h200;
			16'h7f6d: y = 16'h200;
			16'h7f6e: y = 16'h200;
			16'h7f6f: y = 16'h200;
			16'h7f70: y = 16'h200;
			16'h7f71: y = 16'h200;
			16'h7f72: y = 16'h200;
			16'h7f73: y = 16'h200;
			16'h7f74: y = 16'h200;
			16'h7f75: y = 16'h200;
			16'h7f76: y = 16'h200;
			16'h7f77: y = 16'h200;
			16'h7f78: y = 16'h200;
			16'h7f79: y = 16'h200;
			16'h7f7a: y = 16'h200;
			16'h7f7b: y = 16'h200;
			16'h7f7c: y = 16'h200;
			16'h7f7d: y = 16'h200;
			16'h7f7e: y = 16'h200;
			16'h7f7f: y = 16'h200;
			16'h7f80: y = 16'h200;
			16'h7f81: y = 16'h200;
			16'h7f82: y = 16'h200;
			16'h7f83: y = 16'h200;
			16'h7f84: y = 16'h200;
			16'h7f85: y = 16'h200;
			16'h7f86: y = 16'h200;
			16'h7f87: y = 16'h200;
			16'h7f88: y = 16'h200;
			16'h7f89: y = 16'h200;
			16'h7f8a: y = 16'h200;
			16'h7f8b: y = 16'h200;
			16'h7f8c: y = 16'h200;
			16'h7f8d: y = 16'h200;
			16'h7f8e: y = 16'h200;
			16'h7f8f: y = 16'h200;
			16'h7f90: y = 16'h200;
			16'h7f91: y = 16'h200;
			16'h7f92: y = 16'h200;
			16'h7f93: y = 16'h200;
			16'h7f94: y = 16'h200;
			16'h7f95: y = 16'h200;
			16'h7f96: y = 16'h200;
			16'h7f97: y = 16'h200;
			16'h7f98: y = 16'h200;
			16'h7f99: y = 16'h200;
			16'h7f9a: y = 16'h200;
			16'h7f9b: y = 16'h200;
			16'h7f9c: y = 16'h200;
			16'h7f9d: y = 16'h200;
			16'h7f9e: y = 16'h200;
			16'h7f9f: y = 16'h200;
			16'h7fa0: y = 16'h200;
			16'h7fa1: y = 16'h200;
			16'h7fa2: y = 16'h200;
			16'h7fa3: y = 16'h200;
			16'h7fa4: y = 16'h200;
			16'h7fa5: y = 16'h200;
			16'h7fa6: y = 16'h200;
			16'h7fa7: y = 16'h200;
			16'h7fa8: y = 16'h200;
			16'h7fa9: y = 16'h200;
			16'h7faa: y = 16'h200;
			16'h7fab: y = 16'h200;
			16'h7fac: y = 16'h200;
			16'h7fad: y = 16'h200;
			16'h7fae: y = 16'h200;
			16'h7faf: y = 16'h200;
			16'h7fb0: y = 16'h200;
			16'h7fb1: y = 16'h200;
			16'h7fb2: y = 16'h200;
			16'h7fb3: y = 16'h200;
			16'h7fb4: y = 16'h200;
			16'h7fb5: y = 16'h200;
			16'h7fb6: y = 16'h200;
			16'h7fb7: y = 16'h200;
			16'h7fb8: y = 16'h200;
			16'h7fb9: y = 16'h200;
			16'h7fba: y = 16'h200;
			16'h7fbb: y = 16'h200;
			16'h7fbc: y = 16'h200;
			16'h7fbd: y = 16'h200;
			16'h7fbe: y = 16'h200;
			16'h7fbf: y = 16'h200;
			16'h7fc0: y = 16'h200;
			16'h7fc1: y = 16'h200;
			16'h7fc2: y = 16'h200;
			16'h7fc3: y = 16'h200;
			16'h7fc4: y = 16'h200;
			16'h7fc5: y = 16'h200;
			16'h7fc6: y = 16'h200;
			16'h7fc7: y = 16'h200;
			16'h7fc8: y = 16'h200;
			16'h7fc9: y = 16'h200;
			16'h7fca: y = 16'h200;
			16'h7fcb: y = 16'h200;
			16'h7fcc: y = 16'h200;
			16'h7fcd: y = 16'h200;
			16'h7fce: y = 16'h200;
			16'h7fcf: y = 16'h200;
			16'h7fd0: y = 16'h200;
			16'h7fd1: y = 16'h200;
			16'h7fd2: y = 16'h200;
			16'h7fd3: y = 16'h200;
			16'h7fd4: y = 16'h200;
			16'h7fd5: y = 16'h200;
			16'h7fd6: y = 16'h200;
			16'h7fd7: y = 16'h200;
			16'h7fd8: y = 16'h200;
			16'h7fd9: y = 16'h200;
			16'h7fda: y = 16'h200;
			16'h7fdb: y = 16'h200;
			16'h7fdc: y = 16'h200;
			16'h7fdd: y = 16'h200;
			16'h7fde: y = 16'h200;
			16'h7fdf: y = 16'h200;
			16'h7fe0: y = 16'h200;
			16'h7fe1: y = 16'h200;
			16'h7fe2: y = 16'h200;
			16'h7fe3: y = 16'h200;
			16'h7fe4: y = 16'h200;
			16'h7fe5: y = 16'h200;
			16'h7fe6: y = 16'h200;
			16'h7fe7: y = 16'h200;
			16'h7fe8: y = 16'h200;
			16'h7fe9: y = 16'h200;
			16'h7fea: y = 16'h200;
			16'h7feb: y = 16'h200;
			16'h7fec: y = 16'h200;
			16'h7fed: y = 16'h200;
			16'h7fee: y = 16'h200;
			16'h7fef: y = 16'h200;
			16'h7ff0: y = 16'h200;
			16'h7ff1: y = 16'h200;
			16'h7ff2: y = 16'h200;
			16'h7ff3: y = 16'h200;
			16'h7ff4: y = 16'h200;
			16'h7ff5: y = 16'h200;
			16'h7ff6: y = 16'h200;
			16'h7ff7: y = 16'h200;
			16'h7ff8: y = 16'h200;
			16'h7ff9: y = 16'h200;
			16'h7ffa: y = 16'h200;
			16'h7ffb: y = 16'h200;
			16'h7ffc: y = 16'h200;
			16'h7ffd: y = 16'h200;
			16'h7ffe: y = 16'h200;
			16'h7fff: y = 16'h200;
			default: y = 0;
		endcase
	end
endmodule
